`timescale  1ns/1ns
//=================================================================================
//  Author       ：la
//  Project name ：Gas Sensor on FPGA
//  Module Name  : tft_pic
//  Created Time ：2022.5.12
//  Description  ：文字和图像生成模块
//=================================================================================

module  tft_pic
(
    input   wire             tft_clk_33m  ,               //输入工作时钟,频率33MHz
    input   wire             sys_rst_n    ,               //输入复位信号,低电平有效
    input   wire    [10:0]   pix_x        ,               //输入TFT有效显示区域像素点X轴坐标
    input   wire    [10:0]   pix_y        ,               //输入TFT有效显示区域像素点Y轴坐标

    input   wire    [9:0]    ch1          ,               //AD数据
    input   wire    [3:0]    unit1        ,               //个位BCD码
    input   wire    [3:0]    ten1         ,               //十位BCD码
    input   wire    [3:0]    hun1         ,               //百位BCD码

    input   wire    [9:0]    ch2          ,               //AD数据
    input   wire    [3:0]    unit2        ,               //个位BCD码
    input   wire    [3:0]    ten2         ,               //十位BCD码
    input   wire    [3:0]    hun2         ,               //百位BCD码  

    input   wire    [9:0]    ch3          ,               //AD数据
    input   wire    [3:0]    unit3        ,               //个位BCD码
    input   wire    [3:0]    ten3         ,               //十位BCD码
    input   wire    [3:0]    hun3         ,               //百位BCD码

    input   wire    [9:0]    ch4          ,               //AD数据
    input   wire    [3:0]    unit4        ,               //个位BCD码
    input   wire    [3:0]    ten4         ,               //十位BCD码
    input   wire    [3:0]    hun4         ,               //百位BCD码   

    input   wire    [3:0]    unit5        ,               //个位BCD码
    input   wire    [3:0]    ten5         ,               //十位BCD码
    input   wire    [3:0]    hun5         ,               //百位BCD码    

    input   wire   [9:0]   data_out       ,            //输出数据给lcd显示
    input   wire   [2:0]   data_flag      ,



    output  reg     [23:0]   pix_data                     //输出像素点色彩信息
);          

//--------------------------------------------------------------------------
//------------------------------参数和变量定义-------------------------------
//--------------------------------------------------------------------------

parameter   H_VALID =   11'd800            ,              //行有效数据
            V_VALID =   11'd480            ;              //场有效数据
//224*24                       
// parameter   CHAR_x1=   10'd296             ,              //JLU GAS SENSOR 开始X轴坐标
//             CHAR_y1=   10'd8               ;              //JLU GAS SENSOR 开始Y轴坐标
//800*24                       
parameter   CHAR_x3=   10'd10               ,              //CH开始X轴坐标
            CHAR_y3=   10'd416             ;              //CH开始Y轴坐标  
//800*24                       
parameter   CHAR_x4=   10'd0               ,              //NH3开始X轴坐标
            CHAR_y4=   10'd448             ;              //NH3开始Y轴坐标  
                 
parameter   BLACK   =  24'h000000          ,              //黑色
            GOLDEN  =  24'h00ffff          ,              //金色
            WHITE   =  24'hffffff          ,              //白色 
            RED     =  24'hff0000          ,
            BLUE     = 24'h0000ff          ;

// parameter WHITE_R       = 8'hff;
// parameter WHITE_G       = 8'hff;
// parameter WHITE_B       = 8'hff;
// parameter YELLOW_R      = 8'hff;
// parameter YELLOW_G      = 8'hff;
// parameter YELLOW_B      = 8'h00;                                
// parameter CYAN_R        = 8'h00;
// parameter CYAN_G        = 8'hff;
// parameter CYAN_B        = 8'hff;                                
// parameter GREEN_R       = 8'h00;
// parameter GREEN_G       = 8'hff;
// parameter GREEN_B       = 8'h00;
// parameter MAGENTA_R     = 8'hff;
// parameter MAGENTA_G     = 8'h00;
// parameter MAGENTA_B     = 8'hff;
// parameter RED_R         = 8'hff;
// parameter RED_G         = 8'h00;
// parameter RED_B         = 8'h00;
// parameter BLUE_R        = 8'h00;
// parameter BLUE_G        = 8'h00;
// parameter BLUE_B        = 8'hff;
// parameter BLACK_R       = 8'h00;
// parameter BLACK_G       = 8'h00;
// parameter BLACK_B       = 8'h00; 
 
wire    [10:0]   char1_x                   ;              //JLU GAS SENSOR显示X轴坐标
wire    [10:0]   char1_y                   ;              //JLU GAS SENSOR显示Y轴坐标
wire    [10:0]   char3_x                   ;              //CH显示X轴坐标
wire    [10:0]   char3_y                   ;              //CH显示Y轴坐标
wire    [10:0]   char4_x                   ;              //NH3显示X轴坐标
wire    [10:0]   char4_y                   ;             
 
wire    [10:0]   char5_x                   ;
wire    [10:0]   char5_y                   ;
wire    [10:0]   char6_x                   ;
wire    [10:0]   char6_y                   ;
wire    [10:0]   char7_x                   ;
wire    [10:0]   char7_y                   ;
wire    [10:0]   char8_x                   ;
wire    [10:0]   char8_y                   ;
wire    [10:0]   char9_x                   ;
wire    [10:0]   char9_y                   ;
wire    [10:0]   char10_x                  ;
wire    [10:0]   char10_y                  ;
wire    [10:0]   char11_x                  ;
wire    [10:0]   char11_y                  ;
wire    [10:0]   char12_x                  ;
wire    [10:0]   char12_y                  ;
wire    [10:0]   char13_x                  ;
wire    [10:0]   char13_y                  ;
wire    [10:0]   char14_x                  ;
wire    [10:0]   char14_y                  ;
wire    [10:0]   char15_x                  ;
wire    [10:0]   char15_y                  ;
wire    [10:0]   char16_x                  ;
wire    [10:0]   char16_y                  ;
wire    [10:0]   char17_x                  ;
wire    [10:0]   char17_y                  ;
wire    [10:0]   char18_x                  ;
wire    [10:0]   char18_y                  ;
wire    [10:0]   char19_x                  ;
wire    [10:0]   char19_y                  ;
wire    [10:0]   char20_x                  ;
wire    [10:0]   char20_y                  ;
wire    [10:0]   char21_x                  ;
wire    [10:0]   char21_y                  ;
wire    [10:0]   char22_x                  ;
wire    [10:0]   char22_y                  ;
wire    [10:0]   char23_x                  ;
wire    [10:0]   char23_y                  ;
wire    [10:0]   char24_x                  ;
wire    [10:0]   char24_y                  ;
wire    [10:0]   char25_x                  ;
wire    [10:0]   char25_y                  ;
wire    [10:0]   char26_x                  ;
wire    [10:0]   char26_y                  ;


 reg     [223:0] char1     [23:0]          ;              //JLU GAS SENSOR数据
 reg     [63:0]  char3     [23:0]          ;              //CH1
 reg     [63:0]  char19    [23:0]          ;              //CH2
 reg     [63:0]  char20    [23:0]          ;              //CH3
 reg     [63:0]  char21    [23:0]          ;              //CH4
 reg     [63:0]  char4     [23:0]          ;              //NH3数据
 reg     [15:0]  char5     [23:0]          ;              //CH1百位
 reg     [15:0]  char6     [23:0]          ;              //CH1十位
 reg     [15:0]  char7     [23:0]          ;              //CH1个位
 reg     [799:0] char8     [359:0]         ;              //AD图像
 reg     [15:0]  char10    [23:0]          ;              //CH2百位
 reg     [15:0]  char11    [23:0]          ;              //CH2十位
 reg     [15:0]  char12    [23:0]          ;              //CH2个位
 reg     [15:0]  char13    [23:0]          ;              //CH3百位
 reg     [15:0]  char14    [23:0]          ;              //CH3十位
 reg     [15:0]  char15    [23:0]          ;              //CH3个位
 reg     [15:0]  char16    [23:0]          ;              //CH4百位
 reg     [15:0]  char17    [23:0]          ;              //CH4十位
 reg     [15:0]  char18    [23:0]          ;              //CH4个位

 reg     [15:0]  char24    [23:0]          ;              //ppm百位
 reg     [15:0]  char25    [23:0]          ;              //ppm十位
 reg     [15:0]  char26    [23:0]          ;              //ppm个位


//  reg     [31:0]  char22    [23:0]          ;              //欧姆个位
 reg     [47:0]  char23    [23:0]          ;              //ppm  

//--------------------------------------------------------------------------
//---------------------------------Main Code--------------------------------
//--------------------------------------------------------------------------

//---------------------------------------------------------------------------
//---------------------------JLU GAS SNESOR显示坐标---------------------------
//---------------------------------------------------------------------------
// assign  char1_x  =   (((pix_x >= CHAR_x1) && (pix_x < (CHAR_x1 + 10'd224)))
//                     && ((pix_y >= CHAR_y1) && (pix_y < (CHAR_y1 + 10'd24))))
//                     ? (pix_x - CHAR_x1) : 11'h3FF;
// assign  char1_y  =   (((pix_x >= CHAR_x1) && (pix_x < (CHAR_x1 + 10'd224)))
//                     && ((pix_y >= CHAR_y1) && (pix_y < (CHAR_y1 + 10'd24))))
//                     ? (pix_y - CHAR_y1) : 11'h3FF;

// //char:JLU GAS SNESOR
// always@(posedge tft_clk_33m)
//     begin
//         char1[0]     <=  224'h00000000000000000000000000000000000000000000000000000000;
//         char1[1]     <=  224'h00000000000000000000000000000000000000000000000000000000;
//         char1[2]     <=  224'h00000000000000000000000000000000000000000000000000000000;
//         char1[3]     <=  224'h00000000000000000000000000000000000000000000000000000000;
//         char1[4]     <=  224'h0FFF00000000000001EC00C007E0000007E00000000007E003E00000;
//         char1[5]     <=  224'h07FF3E007C0E00000F3C01C01C3C00001C3C3FFE7C0F1C3C0E383FFC;
//         char1[6]     <=  224'h00F81C00380C00001C1C03C0381C0000381C1C063C06381C1C1C1C1E;
//         char1[7]     <=  224'h00F81C00380C0000380C03E0300C0000300C1C033E06300C380E1C0E;
//         char1[8]     <=  224'h00F81C00380C0000380603E03000000030001C0037063000380E1C0E;
//         char1[9]     <=  224'h00F81C00380C0000700006603800000038001C1837863800380F1C0E;
//         char1[10]    <=  224'h00F81C00380C0000700006703C0000003C001C1833863C0078071C1C;
//         char1[11]    <=  224'h00F81C00380C0000700006700F8000000F801C3831C60F8078071C38;
//         char1[12]    <=  224'h00F81C00380C000070000C7003F0000003F01FF831E603F078071FE0;
//         char1[13]    <=  224'h00F81C00380C000070300C38007C0000007C1C1830E6007C78071CE0;
//         char1[14]    <=  224'h00F81C00380C0000701E0FF8001C0000001C1C183076001C78071C70;
//         char1[15]    <=  224'h00F81C00380C0000701C1838000E0000000E1C00307E000E38071C70;
//         char1[16]    <=  224'h00F81C00380C0000381C181C600E0000600E1C00303E600E380E1C38;
//         char1[17]    <=  224'h00F81C03380C0000381C181C300E0000300E1C03301E300E380E1C38;
//         char1[18]    <=  224'h00F81C071C0C00001C1C301C380C0000380C1C06301E380C1C0C1C1C;
//         char1[19]    <=  224'h00F81C0E1C3800000E1C301E3C1C00003C1C1C0E300E3C1C0E381C1C;
//         char1[20]    <=  224'h78F87FFE07E0000003F0FC3F37F0000037F07FFEFC0637F003E07F0F;
//         char1[21]    <=  224'hFCF00000000000000000000000000000000000000000000000000000;
//         char1[22]    <=  224'h7FE00000000000000000000000000000000000000000000000000000;
//         char1[23]    <=  224'h3F800000000000000000000000000000000000000000000000000000;

//     end
//----------------------------------------------------------------------------
//-------------------------------------标尺-----------------------------------
//----------------------------------------------------------------------------
wire    [10:0]   char27_x                  ;
wire    [10:0]   char27_y                  ;
wire    [10:0]   char28_x                  ;
wire    [10:0]   char28_y                  ;
wire    [10:0]   char29_x                  ;
wire    [10:0]   char29_y                  ;
wire    [10:0]   char30_x                  ;
wire    [10:0]   char30_y                  ;
wire    [10:0]   char31_x                  ;
wire    [10:0]   char31_y                  ;
wire    [10:0]   char32_x                  ;
wire    [10:0]   char32_y                  ;

reg     [47:0]  char27    [23:0]          ;              
reg     [47:0]  char28    [23:0]          ;              
reg     [47:0]  char29    [23:0]          ;
reg     [15:0]  char30    [23:0]          ;              
reg     [95:0]  char31    [23:0]          ;              
reg     [95:0]  char32    [23:0]          ;






//char:300
assign  char27_x  =   (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd71) && (pix_y < 10'd95)))
                    ? (pix_x) : 11'h3FF;
assign  char27_y  =    (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd71) && (pix_y < 10'd95)))
                    ? (pix_y - 10'd71) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char27[0]     <=48'h000000000000;
        char27[1]     <=48'h000000000000;
        char27[2]     <=48'h000000000000;
        char27[3]     <=48'h000000000000;
        char27[4]     <=48'h07E001800180;
        char27[5]     <=48'h1EF006600660;
        char27[6]     <=48'h38381C181C18;
        char27[7]     <=48'h383C18181818;
        char27[8]     <=48'h383C300C300C;
        char27[9]     <=48'h003C300C300C;
        char27[10]    <=48'h0078300C300C;
        char27[11]    <=48'h03F0300C300C;
        char27[12]    <=48'h03F0300C300C;
        char27[13]    <=48'h0038300C300C;
        char27[14]    <=48'h001C300C300C;
        char27[15]    <=48'h001E300C300C;
        char27[16]    <=48'h381E300C300C;
        char27[17]    <=48'h781E18181818;
        char27[18]    <=48'h783C18181818;
        char27[19]    <=48'h3C780C300C30;
        char27[20]    <=48'h0FE003C003C0;
        char27[21]    <=48'h000000000000;
        char27[22]    <=48'h000000000000;
        char27[23]    <=48'h000000000000;
    end

//char:200
assign  char28_x  =   (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd171) && (pix_y < 10'd195)))
                    ? (pix_x) : 11'h3FF;
assign  char28_y  =    (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                   && ((pix_y >= 10'd171) && (pix_y < 10'd195)))
                   ? (pix_y - 10'd171) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char28[0]     <=48'h000000000000;
        char28[1]     <=48'h000000000000;
        char28[2]     <=48'h000000000000;
        char28[3]     <=48'h000000000000;
        char28[4]     <=48'h07E001800180;
        char28[5]     <=48'h1EF806600660;
        char28[6]     <=48'h383C1C181C18;
        char28[7]     <=48'h781C18181818;
        char28[8]     <=48'h7C1C300C300C;
        char28[9]     <=48'h381C300C300C;
        char28[10]    <=48'h003C300C300C;
        char28[11]    <=48'h0038300C300C;
        char28[12]    <=48'h0070300C300C;
        char28[13]    <=48'h01E0300C300C;
        char28[14]    <=48'h0380300C300C;
        char28[15]    <=48'h0700300C300C;
        char28[16]    <=48'h0E06300C300C;
        char28[17]    <=48'h1C0E18181818;
        char28[18]    <=48'h301C18181818;
        char28[19]    <=48'h7FFC0C300C30;
        char28[20]    <=48'h7FFC03C003C0;
        char28[21]    <=48'h000000000000;
        char28[22]    <=48'h000000000000;
        char28[23]    <=48'h000000000000;
    end

//char:100
assign  char29_x  =   (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd271) && (pix_y < 10'd295)))
                    ? (pix_x) : 11'h3FF;
assign  char29_y  =    (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd271) && (pix_y < 10'd295)))
                    ? (pix_y - 10'd271) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char29[0]     <=48'h000000000000;
        char29[1]     <=48'h000000000000;
        char29[2]     <=48'h000000000000;
        char29[3]     <=48'h000000000000;
        char29[4]     <=48'h00C001800180;
        char29[5]     <=48'h0FC006600660;
        char29[6]     <=48'h1FC01C181C18;
        char29[7]     <=48'h03C018181818;
        char29[8]     <=48'h03C0300C300C;
        char29[9]     <=48'h03C0300C300C;
        char29[10]    <=48'h03C0300C300C;
        char29[11]    <=48'h03C0300C300C;
        char29[12]    <=48'h03C0300C300C;
        char29[13]    <=48'h03C0300C300C;
        char29[14]    <=48'h03C0300C300C;
        char29[15]    <=48'h03C0300C300C;
        char29[16]    <=48'h03C0300C300C;
        char29[17]    <=48'h03C018181818;
        char29[18]    <=48'h03C018181818;
        char29[19]    <=48'h03E00C300C30;
        char29[20]    <=48'h1FFC03C003C0;
        char29[21]    <=48'h000000000000;
        char29[22]    <=48'h000000000000;
        char29[23]    <=48'h000000000000;
    end

//char:0
assign  char30_x  =   (((pix_x >= 10'd16) && (pix_x < (10'd32)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395)))
                    ? (pix_x-10'd16) : 11'h3FF;
assign  char30_y  =    (((pix_x >= 10'd16) && (pix_x < (10'd32)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395)))
                    ? (pix_y - 10'd371) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char30[0]     <=16'h0000;
        char30[1]     <=16'h0000;
        char30[2]     <=16'h0000;
        char30[3]     <=16'h0000;
        char30[4]     <=16'h07E0;
        char30[5]     <=16'h0FF0;
        char30[6]     <=16'h1C38;
        char30[7]     <=16'h3C3C;
        char30[8]     <=16'h781C;
        char30[9]     <=16'h781E;
        char30[10]    <=16'h781E;
        char30[11]    <=16'h781E;
        char30[12]    <=16'h781E;
        char30[13]    <=16'h781E;
        char30[14]    <=16'h781E;
        char30[15]    <=16'h781E;
        char30[16]    <=16'h781E;
        char30[17]    <=16'h383C;
        char30[18]    <=16'h3C38;
        char30[19]    <=16'h1E78;
        char30[20]    <=16'h07E0;
        char30[21]    <=16'h0000;
        char30[22]    <=16'h0000;
        char30[23]    <=16'h0000;
    end

//char:10min
assign  char31_x  =   (((pix_x >= 10'd352) && (pix_x < (10'd448)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395)))
                    ? (pix_x-10'd352) : 11'h3FF;
assign  char31_y  =    (((pix_x >= 10'd352) && (pix_x < (10'd448)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395)))
                    ? (pix_y - 10'd371) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char31[0]     <=96'h000000000000000000000000;
        char31[1]     <=96'h000000000000000000000000;
        char31[2]     <=96'h000000000000000000000000;
        char31[3]     <=96'h000000000000000000000000;
        char31[4]     <=96'h00C001800000000001800000;
        char31[5]     <=96'h0FC006600000000001C00000;
        char31[6]     <=96'h1FC01C180000000001800000;
        char31[7]     <=96'h03C018180000000000000000;
        char31[8]     <=96'h03C0300C0000000000000000;
        char31[9]     <=96'h03C0300C0000000000000000;
        char31[10]    <=96'h03C0300C0000EF3C1F807BF0;
        char31[11]    <=96'h03C0300C000031C601801C18;
        char31[12]    <=96'h03C0300C0000218601801818;
        char31[13]    <=96'h03C0300C0000218601801818;
        char31[14]    <=96'h03C0300C0000218601801818;
        char31[15]    <=96'h03C0300C0000218601801818;
        char31[16]    <=96'h03C0300C0000218601801818;
        char31[17]    <=96'h03C018180000218601801818;
        char31[18]    <=96'h03C018180000218601801818;
        char31[19]    <=96'h03E00C300000218601801818;
        char31[20]    <=96'h1FFC03C00000FBCF1FF87C3E;
        char31[21]    <=96'h000000000000000000000000;
        char31[22]    <=96'h000000000000000000000000;
        char31[23]    <=96'h000000000000000000000000;
    end

//char:20min
assign  char32_x  =   (((pix_x >= 10'd652) && (pix_x < (10'd748)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395)))
                    ? (pix_x-10'd652) : 11'h3FF;
assign  char32_y  =    (((pix_x >= 10'd652) && (pix_x < (10'd748)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395)))
                    ? (pix_y - 10'd371) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char32[0]     <=96'h000000000000000000000000;
        char32[1]     <=96'h000000000000000000000000;
        char32[2]     <=96'h000000000000000000000000;
        char32[3]     <=96'h000000000000000000000000;
        char32[4]     <=96'h03C001800000000001800000;
        char32[5]     <=96'h0C3006600000000001C00000;
        char32[6]     <=96'h10181C180000000001800000;
        char32[7]     <=96'h300C18180000000000000000;
        char32[8]     <=96'h380C300C0000000000000000;
        char32[9]     <=96'h381C300C0000000000000000;
        char32[10]    <=96'h0018300C0000EF3C1F807BF0;
        char32[11]    <=96'h0030300C000031C601801C18;
        char32[12]    <=96'h0060300C0000218601801818;
        char32[13]    <=96'h00C0300C0000218601801818;
        char32[14]    <=96'h0180300C0000218601801818;
        char32[15]    <=96'h0200300C0000218601801818;
        char32[16]    <=96'h0400300C0000218601801818;
        char32[17]    <=96'h180418180000218601801818;
        char32[18]    <=96'h300C18180000218601801818;
        char32[19]    <=96'h3FF80C300000218601801818;
        char32[20]    <=96'h3FF803C00000FBCF1FF87C3E;
        char32[21]    <=96'h000000000000000000000000;
        char32[22]    <=96'h000000000000000000000000;
        char32[23]    <=96'h000000000000000000000000;
    end
//-----------------------------------------------------------------------------
//-------------------------------------模式4-----------------------------------
//-----------------------------------------------------------------------------
wire    [10:0]   char33_x                  ;
wire    [10:0]   char33_y                  ;
wire    [10:0]   char34_x                  ;
wire    [10:0]   char34_y                  ;
wire    [10:0]   char35_x                  ;
wire    [10:0]   char35_y                  ;
wire    [10:0]   char36_x                  ;
wire    [10:0]   char36_y                  ;

wire    [10:0]   char37_x                  ;
wire    [10:0]   char37_y                  ;
wire    [10:0]   char38_x                  ;
wire    [10:0]   char38_y                  ;
wire    [10:0]   char39_x                  ;
wire    [10:0]   char39_y                  ;
wire    [10:0]   char40_x                  ;
wire    [10:0]   char40_y                  ;

wire    [10:0]   char41_x                  ;
wire    [10:0]   char41_y                  ;
wire    [10:0]   char42_x                  ;
wire    [10:0]   char42_y                  ;
wire    [10:0]   char43_x                  ;
wire    [10:0]   char43_y                  ;
wire    [10:0]   char44_x                  ;
wire    [10:0]   char44_y                  ;

reg     [47:0]  char33    [15:0]          ;     //10min         
reg     [23:0]  char34    [15:0]          ;      //0        
reg     [23:0]  char35    [15:0]          ;      //100   



//char:10min
always@(posedge tft_clk_33m)
    begin
        char33[0]     <=48'h000000000000;
        char33[1]     <=48'h000000000000;
        char33[2]     <=48'h000000000000;
        char33[3]     <=48'h081800003000;
        char33[4]     <=48'h382400003000;
        char33[5]     <=48'h084200000000;
        char33[6]     <=48'h084200000000;
        char33[7]     <=48'h084200FE70DC;
        char33[8]     <=48'h084200491062;
        char33[9]     <=48'h084200491042;
        char33[10]    <=48'h084200491042;
        char33[11]    <=48'h084200491042;
        char33[12]    <=48'h082400491042;
        char33[13]    <=48'h3E1800ED7CE7;
        char33[14]    <=48'h000000000000;
        char33[15]    <=48'h000000000000;
    end

//char:0
always@(posedge tft_clk_33m)
    begin
        char34[0]     <=24'h000000;
        char34[1]     <=24'h000000;
        char34[2]     <=24'h000000;
        char34[3]     <=24'h001800;
        char34[4]     <=24'h002400;
        char34[5]     <=24'h004200;
        char34[6]     <=24'h004200;
        char34[7]     <=24'h004200;
        char34[8]     <=24'h004200;
        char34[9]     <=24'h004200;
        char34[10]    <=24'h004200;
        char34[11]    <=24'h004200;
        char34[12]    <=24'h002400;
        char34[13]    <=24'h001800;
        char34[14]    <=24'h000000;
        char34[15]    <=24'h000000;
    end

//char:100
always@(posedge tft_clk_33m)
    begin
        char35[0]     <=24'h000000;
        char35[1]     <=24'h000000;
        char35[2]     <=24'h000000;
        char35[3]     <=24'h081818;
        char35[4]     <=24'h382424;
        char35[5]     <=24'h084242;
        char35[6]     <=24'h084242;
        char35[7]     <=24'h084242;
        char35[8]     <=24'h084242;
        char35[9]     <=24'h084242;
        char35[10]    <=24'h084242;
        char35[11]    <=24'h084242;
        char35[12]    <=24'h082424;
        char35[13]    <=24'h3E1818;
        char35[14]    <=24'h000000;
        char35[15]    <=24'h000000;
    end

assign  char33_x  =   (((pix_x >= 10'd201) && (pix_x < (10'd249)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_x-10'd201) : 11'h3FF;
assign  char33_y  =    (((pix_x >= 10'd201) && (pix_x < (10'd249)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_y - 10'd165) : 11'h3FF;
assign  char34_x  =   (((pix_x >= 10'd601) && (pix_x < (10'd649)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_x-10'd601) : 11'h3FF;
assign  char34_y  =    (((pix_x >= 10'd601) && (pix_x < (10'd649)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_y - 10'd165) : 11'h3FF;
assign  char35_x  =  (((pix_x >= 10'd201) && (pix_x < (10'd249)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_x-10'd201) : 11'h3FF;
assign  char35_y  =   (((pix_x >= 10'd201) && (pix_x < (10'd249)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_y-10'd345) : 11'h3FF;
assign  char36_x  =   (((pix_x >= 10'd601) && (pix_x < (10'd649)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_x-10'd601) : 11'h3FF;
assign  char36_y  =    (((pix_x >= 10'd601) && (pix_x < (10'd649)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_y - 10'd345) : 11'h3FF;

assign  char37_x  =   (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_x-10'd21) : 11'h3FF;
assign  char37_y  =     (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_y - 10'd165) : 11'h3FF;
assign  char38_x  =   (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_x-10'd421) : 11'h3FF;
assign  char38_y  =   (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))
                    ? (pix_y - 10'd165) : 11'h3FF;
assign  char39_x  =   (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_x-10'd21) : 11'h3FF;
assign  char39_y  =    (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_y - 10'd345) : 11'h3FF;
assign  char40_x  = (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_x-10'd421) : 11'h3FF;
assign  char40_y  =  (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))
                    ? (pix_y - 10'd345) : 11'h3FF;

assign  char41_x  =   (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd115) && (pix_y < 10'd131)))
                    ? (pix_x-10'd21) : 11'h3FF;
assign  char41_y  =   (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd115) && (pix_y < 10'd131)))
                    ? (pix_y - 10'd115) : 11'h3FF;
assign  char42_x  =   (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd115) && (pix_y < 10'd131)))
                    ? (pix_x-10'd421) : 11'h3FF;
assign  char42_y  =   (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd115) && (pix_y < 10'd131)))
                    ? (pix_y - 10'd115) : 11'h3FF;
assign  char43_x  = (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd295) && (pix_y < 10'd311)))
                    ? (pix_x-10'd21) : 11'h3FF;
assign  char43_y  =  (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd295) && (pix_y < 10'd311)))
                    ? (pix_y - 10'd295) : 11'h3FF;
assign  char44_x  =  (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd295) && (pix_y < 10'd311)))
                    ? (pix_x-10'd421) : 11'h3FF;
assign  char44_y  =  (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd295) && (pix_y < 10'd311)))
                    ? (pix_y - 10'd295) : 11'h3FF;

//---------------------------------------------------------------------------
//---------------------------------CH显示坐标---------------------------------
//---------------------------------------------------------------------------

//char:CH1
assign  char3_x  =   (((pix_x >= CHAR_x3) && (pix_x < (10'd74)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_x - CHAR_x3) : 11'h3FF;
assign  char3_y  =   (((pix_x >= CHAR_x3) && (pix_x < (10'd74)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_y - CHAR_y3) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char3[0]     <=64'h0000000000000000;
        char3[1]     <=64'h0000000000000000;
        char3[2]     <=64'h0000000000000000;
        char3[3]     <=64'h0000000000000000;
        char3[4]     <=64'h01E0000000800000;
        char3[5]     <=64'h061C381C01800000;
        char3[6]     <=64'h1804300C07800000;
        char3[7]     <=64'h1806300C01800000;
        char3[8]     <=64'h3002300C01800000;
        char3[9]     <=64'h3000300C01800100;
        char3[10]    <=64'h7000300C01800380;
        char3[11]    <=64'h6000300C01800380;
        char3[12]    <=64'h60003FFC01800000;
        char3[13]    <=64'h6000300C01800000;
        char3[14]    <=64'h6000300C01800000;
        char3[15]    <=64'h7000300C01800000;
        char3[16]    <=64'h3002300C01800000;
        char3[17]    <=64'h3004300C01800000;
        char3[18]    <=64'h1804300C01800180;
        char3[19]    <=64'h0C18300C01C00380;
        char3[20]    <=64'h03E0FC3E0FF80380;
        char3[21]    <=64'h0000000000000000;
        char3[22]    <=64'h0000000000000000;
        char3[23]    <=64'h0000000000000000;
    end

//char:CH2
assign  char19_x  =   (((pix_x >= 10'd200) && (pix_x < (10'd264)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_x - 10'd200) : 11'h3FF;
assign  char19_y  =   (((pix_x >= 10'd200) && (pix_x < (10'd264)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_y - CHAR_y3) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char19[0]     <=64'h0000000000000000;
        char19[1]     <=64'h0000000000000000;
        char19[2]     <=64'h0000000000000000;
        char19[3]     <=64'h0000000000000000;
        char19[4]     <=64'h03FE000003C00000;
        char19[5]     <=64'h0F3E381C0C300000;
        char19[6]     <=64'h1C0E300C10180000;
        char19[7]     <=64'h3806300C300C0000;
        char19[8]     <=64'h7807300C380C0000;
        char19[9]     <=64'h7800300C381C0100;
        char19[10]    <=64'hF000300C00180380;
        char19[11]    <=64'hF000300C00300380;
        char19[12]    <=64'hF0003FFC00600000;
        char19[13]    <=64'hF000300C00C00000;
        char19[14]    <=64'hF000300C01800000;
        char19[15]    <=64'h7000300C02000000;
        char19[16]    <=64'h7807300C04000000;
        char19[17]    <=64'h7806300C18040000;
        char19[18]    <=64'h3C0C300C300C0180;
        char19[19]    <=64'h1F3C300C3FF80380;
        char19[20]    <=64'h07F0FC3E3FF80380;
        char19[21]    <=64'h0000000000000000;
        char19[22]    <=64'h0000000000000000;
        char19[23]    <=64'h0000000000000000;
    end

//char:CH3
assign  char20_x  =   (((pix_x >= 10'd400) && (pix_x < (10'd464)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_x - 10'd400) : 11'h3FF;
assign  char20_y  =   (((pix_x >= 10'd400) && (pix_x < (10'd464)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_y - CHAR_y3) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char20[0]     <=64'h0000000000000000;
        char20[1]     <=64'h0000000000000000;
        char20[2]     <=64'h0000000000000000;
        char20[3]     <=64'h0000000000000000;
        char20[4]     <=64'h03FE000007800000;
        char20[5]     <=64'h0F3E381C08700000;
        char20[6]     <=64'h1C0E300C10380000;
        char20[7]     <=64'h3806300C38180000;
        char20[8]     <=64'h7807300C18180000;
        char20[9]     <=64'h7800300C00180100;
        char20[10]    <=64'hF000300C00300380;
        char20[11]    <=64'hF000300C00E00380;
        char20[12]    <=64'hF0003FFC01E00000;
        char20[13]    <=64'hF000300C00180000;
        char20[14]    <=64'hF000300C00180000;
        char20[15]    <=64'h7000300C000C0000;
        char20[16]    <=64'h7807300C100C0000;
        char20[17]    <=64'h7806300C380C0000;
        char20[18]    <=64'h3C0C300C30180180;
        char20[19]    <=64'h1F3C300C18300380;
        char20[20]    <=64'h07F0FC3E07C00380;
        char20[21]    <=64'h0000000000000000;
        char20[22]    <=64'h0000000000000000;
        char20[23]    <=64'h0000000000000000;
    end

//char:CH4
assign  char21_x  =   (((pix_x >= 10'd600) && (pix_x < (10'd664)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_x - 10'd600) : 11'h3FF;
assign  char21_y  =   (((pix_x >= 10'd600) && (pix_x < (10'd664)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
                    ? (pix_y - CHAR_y3) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char21[0]     <=64'h0000000000000000;
        char21[1]     <=64'h0000000000000000;
        char21[2]     <=64'h0000000000000000;
        char21[3]     <=64'h0000000000000000;
        char21[4]     <=64'h03FE000000300000;
        char21[5]     <=64'h0F3E381C00700000;
        char21[6]     <=64'h1C0E300C00F00000;
        char21[7]     <=64'h3806300C00F00000;
        char21[8]     <=64'h7807300C01700000;
        char21[9]     <=64'h7800300C02700100;
        char21[10]    <=64'hF000300C04700380;
        char21[11]    <=64'hF000300C08700380;
        char21[12]    <=64'hF0003FFC18700000;
        char21[13]    <=64'hF000300C10700000;
        char21[14]    <=64'hF000300C20700000;
        char21[15]    <=64'h7000300C7FFE0000;
        char21[16]    <=64'h7807300C00700000;
        char21[17]    <=64'h7806300C00700000;
        char21[18]    <=64'h3C0C300C00700180;
        char21[19]    <=64'h1F3C300C00700380;
        char21[20]    <=64'h07F0FC3E03FE0380;
        char21[21]    <=64'h0000000000000000;
        char21[22]    <=64'h0000000000000000;
        char21[23]    <=64'h0000000000000000;
    end
// //char:欧姆22
// assign  char22_x  =   (((pix_x >= 10'd600) && (pix_x < (10'd664)))
//                     && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
//                     ? (pix_x - 10'd600) : 11'h3FF;
// assign  char22_y  =   (((pix_x >= 10'd600) && (pix_x < (10'd664)))
//                     && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
//                     ? (pix_y - CHAR_y3) : 11'h3FF;

// always@(posedge tft_clk_33m)
//     begin
//         char22[0]     <=31'h00000000;
//         char22[1]     <=31'h00000000;
//         char22[2]     <=31'h00000000;
//         char22[3]     <=31'h00000000;
//         char22[4]     <=31'h0007E000;
//         char22[5]     <=31'h00181C00;
//         char22[6]     <=31'h00300E00;
//         char22[7]     <=31'h00600700;
//         char22[8]     <=31'h00C00300;
//         char22[9]     <=31'h00C00300;
//         char22[10]    <=31'h00C00300;
//         char22[11]    <=31'h00C00300;
//         char22[12]    <=31'h00C00300;
//         char22[13]    <=31'h00E00700;
//         char22[14]    <=31'h00700E00;
//         char22[15]    <=31'h001C3800;
//         char22[16]    <=31'h00844100;
//         char22[17]    <=31'h00FC7F00;
//         char22[18]    <=31'h00FC7F00;
//         char22[19]    <=31'h00000000;
//         char22[20]    <=31'h00000000;
//         char22[21]    <=31'h00000000;
//         char22[22]    <=31'h00000000;
//         char22[23]    <=31'h00000000;
//     end

//char:ppm23
assign  char23_x  =   (((pix_x >= 10'd122) && (pix_x < (10'd170)))
                    && ((pix_y >= 10'd448) && (pix_y < 10'd472)))
                    ? (pix_x - 10'd122) : 11'h3FF;
assign  char23_y  =   (((pix_x >= 10'd122) && (pix_x < (10'd170)))
                    && ((pix_y >= 10'd448) && (pix_y < 10'd472)))
                    ? (pix_y - 10'd448) : 11'h3FF;

always@(posedge tft_clk_33m)
    begin
        char23[0]     <=48'h000000000000;
        char23[1]     <=48'h000000000000;
        char23[2]     <=48'h000000000000;
        char23[3]     <=48'h000000000000;
        char23[4]     <=48'h000000000000;
        char23[5]     <=48'h000000000000;
        char23[6]     <=48'h000000000000;
        char23[7]     <=48'h000000000000;
        char23[8]     <=48'h000000000000;
        char23[9]     <=48'h000000000000;
        char23[10]    <=48'h7BE07BE0EF3C;
        char23[11]    <=48'h1C181C1831C6;
        char23[12]    <=48'h180C180C2186;
        char23[13]    <=48'h180C180C2186;
        char23[14]    <=48'h180C180C2186;
        char23[15]    <=48'h180C180C2186;
        char23[16]    <=48'h180C180C2186;
        char23[17]    <=48'h180C180C2186;
        char23[18]    <=48'h180C180C2186;
        char23[19]    <=48'h1C381C382186;
        char23[20]    <=48'h1BC01BC0FBCF;
        char23[21]    <=48'h180018000000;
        char23[22]    <=48'h180018000000;
        char23[23]    <=48'h3C003C000000;
    end
//----------------------------------------------------------------------------
//---------------------------------NH3显示坐标---------------------------------
//----------------------------------------------------------------------------

assign  char4_x  =   (((pix_x >= 10'd10) && (pix_x < 10'd74))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_x-10'd10) : 11'h3FF;
assign  char4_y  =   (((pix_x >= 10'd10) && (pix_x < 10'd74))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_y - CHAR_y4) : 11'h3FF;

//char:NH3
always@(posedge tft_clk_33m)
    begin
        char4[0]     <=  64'h0000000000000000;
        char4[1]     <=  64'h0000000000000000;
        char4[2]     <=  64'h0000000000000000;
        char4[3]     <=  64'h0000000000000000;
        char4[4]     <=  64'h000000001C000000;
        char4[5]     <=  64'h1C0E303063000000;
        char4[6]     <=  64'h0E043030C1800000;
        char4[7]     <=  64'h0E043030C0800000;
        char4[8]     <=  64'h0B043030C0800000;
        char4[9]     <=  64'h0984303001802000;
        char4[10]    <=  64'h0984303001807000;
        char4[11]    <=  64'h08C4303006007000;
        char4[12]    <=  64'h08C43FF00F000000;
        char4[13]    <=  64'h0864303001800000;
        char4[14]    <=  64'h0834303000C00000;
        char4[15]    <=  64'h0834303000C00000;
        char4[16]    <=  64'h081C3030C0C00000;
        char4[17]    <=  64'h081C3030C0C00000;
        char4[18]    <=  64'h080C3030C0C03000;
        char4[19]    <=  64'h0804303041807000;
        char4[20]    <=  64'h3E04F8783E003000;
        char4[21]    <=  64'h0000000000000000;
        char4[22]    <=  64'h0000000000000000;
        char4[23]    <=  64'h0000000000000000;

    end

//---------------------------------------------------------------------------
//-----------------------------------AD数据----------------------------------
//---------------------------------------------------------------------------


//ch1数据
assign  char5_x  =   (((pix_x >= 10'd74) && (pix_x < (10'd90)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd74) : 11'h3FF;
assign  char5_y  =   (((pix_x >= 10'd74) && (pix_x < (10'd90)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char6_x  =   (((pix_x >= 10'd90) && (pix_x < (10'd106)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd90) : 11'h3FF;
assign  char6_y  =   (((pix_x >= 10'd90) && (pix_x < (10'd106)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char7_x  =   (((pix_x >= 10'd106) && (pix_x < (10'd122)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd106) : 11'h3FF;
assign  char7_y  =   (((pix_x >= 10'd106) && (pix_x < (10'd122)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;


//ch2数据
assign  char10_x  =   (((pix_x >= 10'd264) && (pix_x < (10'd280)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd264) : 11'h3FF;
assign  char10_y  =   (((pix_x >= 10'd264) && (pix_x < (10'd280)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char11_x  =   (((pix_x >= 10'd280) && (pix_x < (10'd296)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd280) : 11'h3FF;
assign  char11_y  =   (((pix_x >= 10'd280) && (pix_x < (10'd296)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char12_x  =   (((pix_x >= 10'd296) && (pix_x < (10'd312)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd296) : 11'h3FF;
assign  char12_y  =   (((pix_x >= 10'd296) && (pix_x < (10'd312)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

//ch3数据
assign  char13_x  =   (((pix_x >= 10'd464) && (pix_x < (10'd480)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd464) : 11'h3FF;
assign  char13_y  =   (((pix_x >= 10'd464) && (pix_x < (10'd480)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char14_x  =   (((pix_x >= 10'd480) && (pix_x < (10'd496)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd480) : 11'h3FF;
assign  char14_y  =   (((pix_x >= 10'd480) && (pix_x < (10'd496)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char15_x  =   (((pix_x >= 10'd496) && (pix_x < (10'd512)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd496) : 11'h3FF;
assign  char15_y  =   (((pix_x >= 10'd496) && (pix_x < (10'd512)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

//ch4数据
assign  char16_x  =   (((pix_x >= 10'd664) && (pix_x < (10'd680)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd664) : 11'h3FF;
assign  char16_y  =   (((pix_x >= 10'd664) && (pix_x < (10'd680)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char17_x  =   (((pix_x >= 10'd680) && (pix_x < (10'd696)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd680) : 11'h3FF;
assign  char17_y  =   (((pix_x >= 10'd680) && (pix_x < (10'd696)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

assign  char18_x  =   (((pix_x >= 10'd696) && (pix_x < (10'd712)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_x - 10'd696) : 11'h3FF;
assign  char18_y  =   (((pix_x >= 10'd696) && (pix_x < (10'd712)))
                    && ((pix_y >= 10'd416) && (pix_y < (10'd440))))
                    ? (pix_y - 10'd416) : 11'h3FF;

//ppm数据
assign  char24_x  =   (((pix_x >= 10'd74) && (pix_x < (10'd90)))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_x - 10'd74) : 11'h3FF;
assign  char24_y  =    (((pix_x >= 10'd74) && (pix_x < (10'd90)))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_y - 10'd448) : 11'h3FF;

assign  char25_x  =   (((pix_x >= 10'd90) && (pix_x < (10'd106)))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_x - 10'd90) : 11'h3FF;
assign  char25_y  =   (((pix_x >= 10'd90) && (pix_x < (10'd106)))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_y - 10'd448) : 11'h3FF;

assign  char26_x  =   (((pix_x >= 10'd106) && (pix_x < (10'd122)))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_x - 10'd106) : 11'h3FF;
assign  char26_y  =    (((pix_x >= 10'd106) && (pix_x < (10'd122)))
                    && ((pix_y >= 10'd448) && (pix_y < (10'd472))))
                    ? (pix_y - 10'd448) : 11'h3FF;
//------------------------------------------------------------------------------
//---------------------------------------CH1------------------------------------
//------------------------------------------------------------------------------

always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char5[0]     <=  16'h0000;
       char5[1]     <=  16'h0000;
       char5[2]     <=  16'h0000;
       char5[3]     <=  16'h0000;
       char5[4]     <=  16'h07E0;
       char5[5]     <=  16'h0FF0;
       char5[6]     <=  16'h1C38;
       char5[7]     <=  16'h3C3C;
       char5[8]     <=  16'h781C;
       char5[9]     <=  16'h781E;
       char5[10]    <=  16'h781E;
       char5[11]    <=  16'h781E;
       char5[12]    <=  16'h781E;
       char5[13]    <=  16'h781E;
       char5[14]    <=  16'h781E;
       char5[15]    <=  16'h781E;
       char5[16]    <=  16'h781E;
       char5[17]    <=  16'h383C;
       char5[18]    <=  16'h3C38;
       char5[19]    <=  16'h1E78;
       char5[20]    <=  16'h07E0;
       char5[21]    <=  16'h0000;
       char5[22]    <=  16'h0000;
       char5[23]    <=  16'h0000;
    end
    else    
        case(hun1)
            4'd0  :  begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h07E0;
                char5[5]     <=  16'h0FF0;
                char5[6]     <=  16'h1C38;
                char5[7]     <=  16'h3C3C;
                char5[8]     <=  16'h781C;
                char5[9]     <=  16'h781E;
                char5[10]    <=  16'h781E;
                char5[11]    <=  16'h781E;
                char5[12]    <=  16'h781E;
                char5[13]    <=  16'h781E;
                char5[14]    <=  16'h781E;
                char5[15]    <=  16'h781E;
                char5[16]    <=  16'h781E;
                char5[17]    <=  16'h383C;
                char5[18]    <=  16'h3C38;
                char5[19]    <=  16'h1E78;
                char5[20]    <=  16'h07E0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h00C0;
                char5[5]     <=  16'h0FC0;
                char5[6]     <=  16'h1FC0;
                char5[7]     <=  16'h03C0;
                char5[8]     <=  16'h03C0;
                char5[9]     <=  16'h03C0;
                char5[10]    <=  16'h03C0;
                char5[11]    <=  16'h03C0;
                char5[12]    <=  16'h03C0;
                char5[13]    <=  16'h03C0;
                char5[14]    <=  16'h03C0;
                char5[15]    <=  16'h03C0;
                char5[16]    <=  16'h03C0;
                char5[17]    <=  16'h03C0;
                char5[18]    <=  16'h03C0;
                char5[19]    <=  16'h03E0;
                char5[20]    <=  16'h1FFC;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end
            4'd2  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h07E0;
                char5[5]     <=  16'h1EF8;
                char5[6]     <=  16'h383C;
                char5[7]     <=  16'h781C;
                char5[8]     <=  16'h7C1C;
                char5[9]     <=  16'h381C;
                char5[10]    <=  16'h003C;
                char5[11]    <=  16'h0038;
                char5[12]    <=  16'h0070;
                char5[13]    <=  16'h01E0;
                char5[14]    <=  16'h0380;
                char5[15]    <=  16'h0700;
                char5[16]    <=  16'h0E06;
                char5[17]    <=  16'h1C0E;
                char5[18]    <=  16'h301C;
                char5[19]    <=  16'h7FFC;
                char5[20]    <=  16'h7FFC;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h07E0;
                char5[5]     <=  16'h1EF0;
                char5[6]     <=  16'h3838;
                char5[7]     <=  16'h383C;
                char5[8]     <=  16'h383C;
                char5[9]     <=  16'h003C;
                char5[10]    <=  16'h0078;
                char5[11]    <=  16'h03F0;
                char5[12]    <=  16'h03F0;
                char5[13]    <=  16'h0038;
                char5[14]    <=  16'h001C;
                char5[15]    <=  16'h001E;
                char5[16]    <=  16'h381E;
                char5[17]    <=  16'h781E;
                char5[18]    <=  16'h783C;
                char5[19]    <=  16'h3C78;
                char5[20]    <=  16'h0FE0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h0070;
                char5[5]     <=  16'h0070;
                char5[6]     <=  16'h00F0;
                char5[7]     <=  16'h01F0;
                char5[8]     <=  16'h03F0;
                char5[9]     <=  16'h0770;
                char5[10]    <=  16'h0E70;
                char5[11]    <=  16'h0C70;
                char5[12]    <=  16'h1870;
                char5[13]    <=  16'h3070;
                char5[14]    <=  16'h7070;
                char5[15]    <=  16'hFFFF;
                char5[16]    <=  16'h0070;
                char5[17]    <=  16'h0070;
                char5[18]    <=  16'h0070;
                char5[19]    <=  16'h00F8;
                char5[20]    <=  16'h07FE;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h1FFC;
                char5[5]     <=  16'h1FFC;
                char5[6]     <=  16'h3800;
                char5[7]     <=  16'h3800;
                char5[8]     <=  16'h3800;
                char5[9]     <=  16'h3800;
                char5[10]    <=  16'h3FF0;
                char5[11]    <=  16'h3FF8;
                char5[12]    <=  16'h383C;
                char5[13]    <=  16'h101C;
                char5[14]    <=  16'h001E;
                char5[15]    <=  16'h001E;
                char5[16]    <=  16'h381E;
                char5[17]    <=  16'h781C;
                char5[18]    <=  16'h783C;
                char5[19]    <=  16'h3C78;
                char5[20]    <=  16'h0FF0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h03F0;
                char5[5]     <=  16'h0F38;
                char5[6]     <=  16'h1C3C;
                char5[7]     <=  16'h383C;
                char5[8]     <=  16'h3800;
                char5[9]     <=  16'h7800;
                char5[10]    <=  16'h7BF0;
                char5[11]    <=  16'h7FF8;
                char5[12]    <=  16'h7C3C;
                char5[13]    <=  16'h781E;
                char5[14]    <=  16'h781E;
                char5[15]    <=  16'h781E;
                char5[16]    <=  16'h781E;
                char5[17]    <=  16'h381E;
                char5[18]    <=  16'h3C1C;
                char5[19]    <=  16'h1E38;
                char5[20]    <=  16'h07F0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h3FFE;
                char5[5]     <=  16'h3FFE;
                char5[6]     <=  16'h381C;
                char5[7]     <=  16'h7018;
                char5[8]     <=  16'h7030;
                char5[9]     <=  16'h0070;
                char5[10]    <=  16'h00E0;
                char5[11]    <=  16'h00E0;
                char5[12]    <=  16'h01C0;
                char5[13]    <=  16'h01C0;
                char5[14]    <=  16'h0380;
                char5[15]    <=  16'h0380;
                char5[16]    <=  16'h0780;
                char5[17]    <=  16'h0780;
                char5[18]    <=  16'h0780;
                char5[19]    <=  16'h0780;
                char5[20]    <=  16'h0780;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h07E0;
                char5[5]     <=  16'h1E78;
                char5[6]     <=  16'h381C;
                char5[7]     <=  16'h701E;
                char5[8]     <=  16'h701E;
                char5[9]     <=  16'h781C;
                char5[10]    <=  16'h3E3C;
                char5[11]    <=  16'h1FF0;
                char5[12]    <=  16'h1FF0;
                char5[13]    <=  16'h3CF8;
                char5[14]    <=  16'h783C;
                char5[15]    <=  16'h701E;
                char5[16]    <=  16'h701E;
                char5[17]    <=  16'h701E;
                char5[18]    <=  16'h701C;
                char5[19]    <=  16'h3C38;
                char5[20]    <=  16'h0FF0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h0FE0;
                char5[5]     <=  16'h1EF8;
                char5[6]     <=  16'h3838;
                char5[7]     <=  16'h781C;
                char5[8]     <=  16'h701E;
                char5[9]     <=  16'h701E;
                char5[10]    <=  16'h701E;
                char5[11]    <=  16'h781E;
                char5[12]    <=  16'h783E;
                char5[13]    <=  16'h3FFE;
                char5[14]    <=  16'h0FDE;
                char5[15]    <=  16'h001C;
                char5[16]    <=  16'h003C;
                char5[17]    <=  16'h1838;
                char5[18]    <=  16'h3C78;
                char5[19]    <=  16'h3CF0;
                char5[20]    <=  16'h1FC0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end   
            default:begin
                char5[0]     <=  16'h0000;
                char5[1]     <=  16'h0000;
                char5[2]     <=  16'h0000;
                char5[3]     <=  16'h0000;
                char5[4]     <=  16'h07E0;
                char5[5]     <=  16'h0FF0;
                char5[6]     <=  16'h1C38;
                char5[7]     <=  16'h3C3C;
                char5[8]     <=  16'h781C;
                char5[9]     <=  16'h781E;
                char5[10]    <=  16'h781E;
                char5[11]    <=  16'h781E;
                char5[12]    <=  16'h781E;
                char5[13]    <=  16'h781E;
                char5[14]    <=  16'h781E;
                char5[15]    <=  16'h781E;
                char5[16]    <=  16'h781E;
                char5[17]    <=  16'h383C;
                char5[18]    <=  16'h3C38;
                char5[19]    <=  16'h1E78;
                char5[20]    <=  16'h07E0;
                char5[21]    <=  16'h0000;
                char5[22]    <=  16'h0000;
                char5[23]    <=  16'h0000;
            end
        endcase
always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char6[0]     <=  16'h0000;
       char6[1]     <=  16'h0000;
       char6[2]     <=  16'h0000;
       char6[3]     <=  16'h0000;
       char6[4]     <=  16'h07E0;
       char6[5]     <=  16'h0FF0;
       char6[6]     <=  16'h1C38;
       char6[7]     <=  16'h3C3C;
       char6[8]     <=  16'h781C;
       char6[9]     <=  16'h781E;
       char6[10]    <=  16'h781E;
       char6[11]    <=  16'h781E;
       char6[12]    <=  16'h781E;
       char6[13]    <=  16'h781E;
       char6[14]    <=  16'h781E;
       char6[15]    <=  16'h781E;
       char6[16]    <=  16'h781E;
       char6[17]    <=  16'h383C;
       char6[18]    <=  16'h3C38;
       char6[19]    <=  16'h1E78;
       char6[20]    <=  16'h07E0;
       char6[21]    <=  16'h0000;
       char6[22]    <=  16'h0000;
       char6[23]    <=  16'h0000;
    end
    else    
        case(ten1)
            4'd0  :  begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h07E0;
                char6[5]     <=  16'h0FF0;
                char6[6]     <=  16'h1C38;
                char6[7]     <=  16'h3C3C;
                char6[8]     <=  16'h781C;
                char6[9]     <=  16'h781E;
                char6[10]    <=  16'h781E;
                char6[11]    <=  16'h781E;
                char6[12]    <=  16'h781E;
                char6[13]    <=  16'h781E;
                char6[14]    <=  16'h781E;
                char6[15]    <=  16'h781E;
                char6[16]    <=  16'h781E;
                char6[17]    <=  16'h383C;
                char6[18]    <=  16'h3C38;
                char6[19]    <=  16'h1E78;
                char6[20]    <=  16'h07E0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h00C0;
                char6[5]     <=  16'h0FC0;
                char6[6]     <=  16'h1FC0;
                char6[7]     <=  16'h03C0;
                char6[8]     <=  16'h03C0;
                char6[9]     <=  16'h03C0;
                char6[10]    <=  16'h03C0;
                char6[11]    <=  16'h03C0;
                char6[12]    <=  16'h03C0;
                char6[13]    <=  16'h03C0;
                char6[14]    <=  16'h03C0;
                char6[15]    <=  16'h03C0;
                char6[16]    <=  16'h03C0;
                char6[17]    <=  16'h03C0;
                char6[18]    <=  16'h03C0;
                char6[19]    <=  16'h03E0;
                char6[20]    <=  16'h1FFC;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end
            4'd2  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h07E0;
                char6[5]     <=  16'h1EF8;
                char6[6]     <=  16'h383C;
                char6[7]     <=  16'h781C;
                char6[8]     <=  16'h7C1C;
                char6[9]     <=  16'h381C;
                char6[10]    <=  16'h003C;
                char6[11]    <=  16'h0038;
                char6[12]    <=  16'h0070;
                char6[13]    <=  16'h01E0;
                char6[14]    <=  16'h0380;
                char6[15]    <=  16'h0700;
                char6[16]    <=  16'h0E06;
                char6[17]    <=  16'h1C0E;
                char6[18]    <=  16'h301C;
                char6[19]    <=  16'h7FFC;
                char6[20]    <=  16'h7FFC;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h07E0;
                char6[5]     <=  16'h1EF0;
                char6[6]     <=  16'h3838;
                char6[7]     <=  16'h383C;
                char6[8]     <=  16'h383C;
                char6[9]     <=  16'h003C;
                char6[10]    <=  16'h0078;
                char6[11]    <=  16'h03F0;
                char6[12]    <=  16'h03F0;
                char6[13]    <=  16'h0038;
                char6[14]    <=  16'h001C;
                char6[15]    <=  16'h001E;
                char6[16]    <=  16'h381E;
                char6[17]    <=  16'h781E;
                char6[18]    <=  16'h783C;
                char6[19]    <=  16'h3C78;
                char6[20]    <=  16'h0FE0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h0070;
                char6[5]     <=  16'h0070;
                char6[6]     <=  16'h00F0;
                char6[7]     <=  16'h01F0;
                char6[8]     <=  16'h03F0;
                char6[9]     <=  16'h0770;
                char6[10]    <=  16'h0E70;
                char6[11]    <=  16'h0C70;
                char6[12]    <=  16'h1870;
                char6[13]    <=  16'h3070;
                char6[14]    <=  16'h7070;
                char6[15]    <=  16'hFFFF;
                char6[16]    <=  16'h0070;
                char6[17]    <=  16'h0070;
                char6[18]    <=  16'h0070;
                char6[19]    <=  16'h00F8;
                char6[20]    <=  16'h07FE;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h1FFC;
                char6[5]     <=  16'h1FFC;
                char6[6]     <=  16'h3800;
                char6[7]     <=  16'h3800;
                char6[8]     <=  16'h3800;
                char6[9]     <=  16'h3800;
                char6[10]    <=  16'h3FF0;
                char6[11]    <=  16'h3FF8;
                char6[12]    <=  16'h383C;
                char6[13]    <=  16'h101C;
                char6[14]    <=  16'h001E;
                char6[15]    <=  16'h001E;
                char6[16]    <=  16'h381E;
                char6[17]    <=  16'h781C;
                char6[18]    <=  16'h783C;
                char6[19]    <=  16'h3C78;
                char6[20]    <=  16'h0FF0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h03F0;
                char6[5]     <=  16'h0F38;
                char6[6]     <=  16'h1C3C;
                char6[7]     <=  16'h383C;
                char6[8]     <=  16'h3800;
                char6[9]     <=  16'h7800;
                char6[10]    <=  16'h7BF0;
                char6[11]    <=  16'h7FF8;
                char6[12]    <=  16'h7C3C;
                char6[13]    <=  16'h781E;
                char6[14]    <=  16'h781E;
                char6[15]    <=  16'h781E;
                char6[16]    <=  16'h781E;
                char6[17]    <=  16'h381E;
                char6[18]    <=  16'h3C1C;
                char6[19]    <=  16'h1E38;
                char6[20]    <=  16'h07F0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h3FFE;
                char6[5]     <=  16'h3FFE;
                char6[6]     <=  16'h381C;
                char6[7]     <=  16'h7018;
                char6[8]     <=  16'h7030;
                char6[9]     <=  16'h0070;
                char6[10]    <=  16'h00E0;
                char6[11]    <=  16'h00E0;
                char6[12]    <=  16'h01C0;
                char6[13]    <=  16'h01C0;
                char6[14]    <=  16'h0380;
                char6[15]    <=  16'h0380;
                char6[16]    <=  16'h0780;
                char6[17]    <=  16'h0780;
                char6[18]    <=  16'h0780;
                char6[19]    <=  16'h0780;
                char6[20]    <=  16'h0780;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h07E0;
                char6[5]     <=  16'h1E78;
                char6[6]     <=  16'h381C;
                char6[7]     <=  16'h701E;
                char6[8]     <=  16'h701E;
                char6[9]     <=  16'h781C;
                char6[10]    <=  16'h3E3C;
                char6[11]    <=  16'h1FF0;
                char6[12]    <=  16'h1FF0;
                char6[13]    <=  16'h3CF8;
                char6[14]    <=  16'h783C;
                char6[15]    <=  16'h701E;
                char6[16]    <=  16'h701E;
                char6[17]    <=  16'h701E;
                char6[18]    <=  16'h701C;
                char6[19]    <=  16'h3C38;
                char6[20]    <=  16'h0FF0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h0FE0;
                char6[5]     <=  16'h1EF8;
                char6[6]     <=  16'h3838;
                char6[7]     <=  16'h781C;
                char6[8]     <=  16'h701E;
                char6[9]     <=  16'h701E;
                char6[10]    <=  16'h701E;
                char6[11]    <=  16'h781E;
                char6[12]    <=  16'h783E;
                char6[13]    <=  16'h3FFE;
                char6[14]    <=  16'h0FDE;
                char6[15]    <=  16'h001C;
                char6[16]    <=  16'h003C;
                char6[17]    <=  16'h1838;
                char6[18]    <=  16'h3C78;
                char6[19]    <=  16'h3CF0;
                char6[20]    <=  16'h1FC0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end   
            default:begin
                char6[0]     <=  16'h0000;
                char6[1]     <=  16'h0000;
                char6[2]     <=  16'h0000;
                char6[3]     <=  16'h0000;
                char6[4]     <=  16'h07E0;
                char6[5]     <=  16'h0FF0;
                char6[6]     <=  16'h1C38;
                char6[7]     <=  16'h3C3C;
                char6[8]     <=  16'h781C;
                char6[9]     <=  16'h781E;
                char6[10]    <=  16'h781E;
                char6[11]    <=  16'h781E;
                char6[12]    <=  16'h781E;
                char6[13]    <=  16'h781E;
                char6[14]    <=  16'h781E;
                char6[15]    <=  16'h781E;
                char6[16]    <=  16'h781E;
                char6[17]    <=  16'h383C;
                char6[18]    <=  16'h3C38;
                char6[19]    <=  16'h1E78;
                char6[20]    <=  16'h07E0;
                char6[21]    <=  16'h0000;
                char6[22]    <=  16'h0000;
                char6[23]    <=  16'h0000;
            end
        endcase

always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char7[0]     <=  16'h0000;
       char7[1]     <=  16'h0000;
       char7[2]     <=  16'h0000;
       char7[3]     <=  16'h0000;
       char7[4]     <=  16'h07E0;
       char7[5]     <=  16'h0FF0;
       char7[6]     <=  16'h1C38;
       char7[7]     <=  16'h3C3C;
       char7[8]     <=  16'h781C;
       char7[9]     <=  16'h781E;
       char7[10]    <=  16'h781E;
       char7[11]    <=  16'h781E;
       char7[12]    <=  16'h781E;
       char7[13]    <=  16'h781E;
       char7[14]    <=  16'h781E;
       char7[15]    <=  16'h781E;
       char7[16]    <=  16'h781E;
       char7[17]    <=  16'h383C;
       char7[18]    <=  16'h3C38;
       char7[19]    <=  16'h1E78;
       char7[20]    <=  16'h07E0;
       char7[21]    <=  16'h0000;
       char7[22]    <=  16'h0000;
       char7[23]    <=  16'h0000;
    end
    else    
        case(unit1)
            4'd0  :  begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h07E0;
                char7[5]     <=  16'h0FF0;
                char7[6]     <=  16'h1C38;
                char7[7]     <=  16'h3C3C;
                char7[8]     <=  16'h781C;
                char7[9]     <=  16'h781E;
                char7[10]    <=  16'h781E;
                char7[11]    <=  16'h781E;
                char7[12]    <=  16'h781E;
                char7[13]    <=  16'h781E;
                char7[14]    <=  16'h781E;
                char7[15]    <=  16'h781E;
                char7[16]    <=  16'h781E;
                char7[17]    <=  16'h383C;
                char7[18]    <=  16'h3C38;
                char7[19]    <=  16'h1E78;
                char7[20]    <=  16'h07E0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h00C0;
                char7[5]     <=  16'h0FC0;
                char7[6]     <=  16'h1FC0;
                char7[7]     <=  16'h03C0;
                char7[8]     <=  16'h03C0;
                char7[9]     <=  16'h03C0;
                char7[10]    <=  16'h03C0;
                char7[11]    <=  16'h03C0;
                char7[12]    <=  16'h03C0;
                char7[13]    <=  16'h03C0;
                char7[14]    <=  16'h03C0;
                char7[15]    <=  16'h03C0;
                char7[16]    <=  16'h03C0;
                char7[17]    <=  16'h03C0;
                char7[18]    <=  16'h03C0;
                char7[19]    <=  16'h03E0;
                char7[20]    <=  16'h1FFC;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end
            4'd2  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h07E0;
                char7[5]     <=  16'h1EF8;
                char7[6]     <=  16'h383C;
                char7[7]     <=  16'h781C;
                char7[8]     <=  16'h7C1C;
                char7[9]     <=  16'h381C;
                char7[10]    <=  16'h003C;
                char7[11]    <=  16'h0038;
                char7[12]    <=  16'h0070;
                char7[13]    <=  16'h01E0;
                char7[14]    <=  16'h0380;
                char7[15]    <=  16'h0700;
                char7[16]    <=  16'h0E06;
                char7[17]    <=  16'h1C0E;
                char7[18]    <=  16'h301C;
                char7[19]    <=  16'h7FFC;
                char7[20]    <=  16'h7FFC;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h07E0;
                char7[5]     <=  16'h1EF0;
                char7[6]     <=  16'h3838;
                char7[7]     <=  16'h383C;
                char7[8]     <=  16'h383C;
                char7[9]     <=  16'h003C;
                char7[10]    <=  16'h0078;
                char7[11]    <=  16'h03F0;
                char7[12]    <=  16'h03F0;
                char7[13]    <=  16'h0038;
                char7[14]    <=  16'h001C;
                char7[15]    <=  16'h001E;
                char7[16]    <=  16'h381E;
                char7[17]    <=  16'h781E;
                char7[18]    <=  16'h783C;
                char7[19]    <=  16'h3C78;
                char7[20]    <=  16'h0FE0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h0070;
                char7[5]     <=  16'h0070;
                char7[6]     <=  16'h00F0;
                char7[7]     <=  16'h01F0;
                char7[8]     <=  16'h03F0;
                char7[9]     <=  16'h0770;
                char7[10]    <=  16'h0E70;
                char7[11]    <=  16'h0C70;
                char7[12]    <=  16'h1870;
                char7[13]    <=  16'h3070;
                char7[14]    <=  16'h7070;
                char7[15]    <=  16'hFFFF;
                char7[16]    <=  16'h0070;
                char7[17]    <=  16'h0070;
                char7[18]    <=  16'h0070;
                char7[19]    <=  16'h00F8;
                char7[20]    <=  16'h07FE;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h1FFC;
                char7[5]     <=  16'h1FFC;
                char7[6]     <=  16'h3800;
                char7[7]     <=  16'h3800;
                char7[8]     <=  16'h3800;
                char7[9]     <=  16'h3800;
                char7[10]    <=  16'h3FF0;
                char7[11]    <=  16'h3FF8;
                char7[12]    <=  16'h383C;
                char7[13]    <=  16'h101C;
                char7[14]    <=  16'h001E;
                char7[15]    <=  16'h001E;
                char7[16]    <=  16'h381E;
                char7[17]    <=  16'h781C;
                char7[18]    <=  16'h783C;
                char7[19]    <=  16'h3C78;
                char7[20]    <=  16'h0FF0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h03F0;
                char7[5]     <=  16'h0F38;
                char7[6]     <=  16'h1C3C;
                char7[7]     <=  16'h383C;
                char7[8]     <=  16'h3800;
                char7[9]     <=  16'h7800;
                char7[10]    <=  16'h7BF0;
                char7[11]    <=  16'h7FF8;
                char7[12]    <=  16'h7C3C;
                char7[13]    <=  16'h781E;
                char7[14]    <=  16'h781E;
                char7[15]    <=  16'h781E;
                char7[16]    <=  16'h781E;
                char7[17]    <=  16'h381E;
                char7[18]    <=  16'h3C1C;
                char7[19]    <=  16'h1E38;
                char7[20]    <=  16'h07F0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h3FFE;
                char7[5]     <=  16'h3FFE;
                char7[6]     <=  16'h381C;
                char7[7]     <=  16'h7018;
                char7[8]     <=  16'h7030;
                char7[9]     <=  16'h0070;
                char7[10]    <=  16'h00E0;
                char7[11]    <=  16'h00E0;
                char7[12]    <=  16'h01C0;
                char7[13]    <=  16'h01C0;
                char7[14]    <=  16'h0380;
                char7[15]    <=  16'h0380;
                char7[16]    <=  16'h0780;
                char7[17]    <=  16'h0780;
                char7[18]    <=  16'h0780;
                char7[19]    <=  16'h0780;
                char7[20]    <=  16'h0780;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h07E0;
                char7[5]     <=  16'h1E78;
                char7[6]     <=  16'h381C;
                char7[7]     <=  16'h701E;
                char7[8]     <=  16'h701E;
                char7[9]     <=  16'h781C;
                char7[10]    <=  16'h3E3C;
                char7[11]    <=  16'h1FF0;
                char7[12]    <=  16'h1FF0;
                char7[13]    <=  16'h3CF8;
                char7[14]    <=  16'h783C;
                char7[15]    <=  16'h701E;
                char7[16]    <=  16'h701E;
                char7[17]    <=  16'h701E;
                char7[18]    <=  16'h701C;
                char7[19]    <=  16'h3C38;
                char7[20]    <=  16'h0FF0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h0FE0;
                char7[5]     <=  16'h1EF8;
                char7[6]     <=  16'h3838;
                char7[7]     <=  16'h781C;
                char7[8]     <=  16'h701E;
                char7[9]     <=  16'h701E;
                char7[10]    <=  16'h701E;
                char7[11]    <=  16'h781E;
                char7[12]    <=  16'h783E;
                char7[13]    <=  16'h3FFE;
                char7[14]    <=  16'h0FDE;
                char7[15]    <=  16'h001C;
                char7[16]    <=  16'h003C;
                char7[17]    <=  16'h1838;
                char7[18]    <=  16'h3C78;
                char7[19]    <=  16'h3CF0;
                char7[20]    <=  16'h1FC0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end   
            default:begin
                char7[0]     <=  16'h0000;
                char7[1]     <=  16'h0000;
                char7[2]     <=  16'h0000;
                char7[3]     <=  16'h0000;
                char7[4]     <=  16'h07E0;
                char7[5]     <=  16'h0FF0;
                char7[6]     <=  16'h1C38;
                char7[7]     <=  16'h3C3C;
                char7[8]     <=  16'h781C;
                char7[9]     <=  16'h781E;
                char7[10]    <=  16'h781E;
                char7[11]    <=  16'h781E;
                char7[12]    <=  16'h781E;
                char7[13]    <=  16'h781E;
                char7[14]    <=  16'h781E;
                char7[15]    <=  16'h781E;
                char7[16]    <=  16'h781E;
                char7[17]    <=  16'h383C;
                char7[18]    <=  16'h3C38;
                char7[19]    <=  16'h1E78;
                char7[20]    <=  16'h07E0;
                char7[21]    <=  16'h0000;
                char7[22]    <=  16'h0000;
                char7[23]    <=  16'h0000;
            end
        endcase

//------------------------------------------------------------------------------
//--------------------------------------CH2-------------------------------------
//------------------------------------------------------------------------------


always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char10[0]     <=  16'h0000;
       char10[1]     <=  16'h0000;
       char10[2]     <=  16'h0000;
       char10[3]     <=  16'h0000;
       char10[4]     <=  16'h07E0;
       char10[5]     <=  16'h0FF0;
       char10[6]     <=  16'h1C38;
       char10[7]     <=  16'h3C3C;
       char10[8]     <=  16'h781C;
       char10[9]     <=  16'h781E;
       char10[10]    <=  16'h781E;
       char10[11]    <=  16'h781E;
       char10[12]    <=  16'h781E;
       char10[13]    <=  16'h781E;
       char10[14]    <=  16'h781E;
       char10[15]    <=  16'h781E;
       char10[16]    <=  16'h781E;
       char10[17]    <=  16'h383C;
       char10[18]    <=  16'h3C38;
       char10[19]    <=  16'h1E78;
       char10[20]    <=  16'h07E0;
       char10[21]    <=  16'h0000;
       char10[22]    <=  16'h0000;
       char10[23]    <=  16'h0000;
    end
    else    
        case(hun2)
            4'd0  :  begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h07E0;
                char10[5]     <=  16'h0FF0;
                char10[6]     <=  16'h1C38;
                char10[7]     <=  16'h3C3C;
                char10[8]     <=  16'h781C;
                char10[9]     <=  16'h781E;
                char10[10]    <=  16'h781E;
                char10[11]    <=  16'h781E;
                char10[12]    <=  16'h781E;
                char10[13]    <=  16'h781E;
                char10[14]    <=  16'h781E;
                char10[15]    <=  16'h781E;
                char10[16]    <=  16'h781E;
                char10[17]    <=  16'h383C;
                char10[18]    <=  16'h3C38;
                char10[19]    <=  16'h1E78;
                char10[20]    <=  16'h07E0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h00C0;
                char10[5]     <=  16'h0FC0;
                char10[6]     <=  16'h1FC0;
                char10[7]     <=  16'h03C0;
                char10[8]     <=  16'h03C0;
                char10[9]     <=  16'h03C0;
                char10[10]    <=  16'h03C0;
                char10[11]    <=  16'h03C0;
                char10[12]    <=  16'h03C0;
                char10[13]    <=  16'h03C0;
                char10[14]    <=  16'h03C0;
                char10[15]    <=  16'h03C0;
                char10[16]    <=  16'h03C0;
                char10[17]    <=  16'h03C0;
                char10[18]    <=  16'h03C0;
                char10[19]    <=  16'h03E0;
                char10[20]    <=  16'h1FFC;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end
            4'd2  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h07E0;
                char10[5]     <=  16'h1EF8;
                char10[6]     <=  16'h383C;
                char10[7]     <=  16'h781C;
                char10[8]     <=  16'h7C1C;
                char10[9]     <=  16'h381C;
                char10[10]    <=  16'h003C;
                char10[11]    <=  16'h0038;
                char10[12]    <=  16'h0070;
                char10[13]    <=  16'h01E0;
                char10[14]    <=  16'h0380;
                char10[15]    <=  16'h0700;
                char10[16]    <=  16'h0E06;
                char10[17]    <=  16'h1C0E;
                char10[18]    <=  16'h301C;
                char10[19]    <=  16'h7FFC;
                char10[20]    <=  16'h7FFC;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h07E0;
                char10[5]     <=  16'h1EF0;
                char10[6]     <=  16'h3838;
                char10[7]     <=  16'h383C;
                char10[8]     <=  16'h383C;
                char10[9]     <=  16'h003C;
                char10[10]    <=  16'h0078;
                char10[11]    <=  16'h03F0;
                char10[12]    <=  16'h03F0;
                char10[13]    <=  16'h0038;
                char10[14]    <=  16'h001C;
                char10[15]    <=  16'h001E;
                char10[16]    <=  16'h381E;
                char10[17]    <=  16'h781E;
                char10[18]    <=  16'h783C;
                char10[19]    <=  16'h3C78;
                char10[20]    <=  16'h0FE0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h0070;
                char10[5]     <=  16'h0070;
                char10[6]     <=  16'h00F0;
                char10[7]     <=  16'h01F0;
                char10[8]     <=  16'h03F0;
                char10[9]     <=  16'h0770;
                char10[10]    <=  16'h0E70;
                char10[11]    <=  16'h0C70;
                char10[12]    <=  16'h1870;
                char10[13]    <=  16'h3070;
                char10[14]    <=  16'h7070;
                char10[15]    <=  16'hFFFF;
                char10[16]    <=  16'h0070;
                char10[17]    <=  16'h0070;
                char10[18]    <=  16'h0070;
                char10[19]    <=  16'h00F8;
                char10[20]    <=  16'h07FE;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h1FFC;
                char10[5]     <=  16'h1FFC;
                char10[6]     <=  16'h3800;
                char10[7]     <=  16'h3800;
                char10[8]     <=  16'h3800;
                char10[9]     <=  16'h3800;
                char10[10]    <=  16'h3FF0;
                char10[11]    <=  16'h3FF8;
                char10[12]    <=  16'h383C;
                char10[13]    <=  16'h101C;
                char10[14]    <=  16'h001E;
                char10[15]    <=  16'h001E;
                char10[16]    <=  16'h381E;
                char10[17]    <=  16'h781C;
                char10[18]    <=  16'h783C;
                char10[19]    <=  16'h3C78;
                char10[20]    <=  16'h0FF0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h03F0;
                char10[5]     <=  16'h0F38;
                char10[6]     <=  16'h1C3C;
                char10[7]     <=  16'h383C;
                char10[8]     <=  16'h3800;
                char10[9]     <=  16'h7800;
                char10[10]    <=  16'h7BF0;
                char10[11]    <=  16'h7FF8;
                char10[12]    <=  16'h7C3C;
                char10[13]    <=  16'h781E;
                char10[14]    <=  16'h781E;
                char10[15]    <=  16'h781E;
                char10[16]    <=  16'h781E;
                char10[17]    <=  16'h381E;
                char10[18]    <=  16'h3C1C;
                char10[19]    <=  16'h1E38;
                char10[20]    <=  16'h07F0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h3FFE;
                char10[5]     <=  16'h3FFE;
                char10[6]     <=  16'h381C;
                char10[7]     <=  16'h7018;
                char10[8]     <=  16'h7030;
                char10[9]     <=  16'h0070;
                char10[10]    <=  16'h00E0;
                char10[11]    <=  16'h00E0;
                char10[12]    <=  16'h01C0;
                char10[13]    <=  16'h01C0;
                char10[14]    <=  16'h0380;
                char10[15]    <=  16'h0380;
                char10[16]    <=  16'h0780;
                char10[17]    <=  16'h0780;
                char10[18]    <=  16'h0780;
                char10[19]    <=  16'h0780;
                char10[20]    <=  16'h0780;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h07E0;
                char10[5]     <=  16'h1E78;
                char10[6]     <=  16'h381C;
                char10[7]     <=  16'h701E;
                char10[8]     <=  16'h701E;
                char10[9]     <=  16'h781C;
                char10[10]    <=  16'h3E3C;
                char10[11]    <=  16'h1FF0;
                char10[12]    <=  16'h1FF0;
                char10[13]    <=  16'h3CF8;
                char10[14]    <=  16'h783C;
                char10[15]    <=  16'h701E;
                char10[16]    <=  16'h701E;
                char10[17]    <=  16'h701E;
                char10[18]    <=  16'h701C;
                char10[19]    <=  16'h3C38;
                char10[20]    <=  16'h0FF0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h0FE0;
                char10[5]     <=  16'h1EF8;
                char10[6]     <=  16'h3838;
                char10[7]     <=  16'h781C;
                char10[8]     <=  16'h701E;
                char10[9]     <=  16'h701E;
                char10[10]    <=  16'h701E;
                char10[11]    <=  16'h781E;
                char10[12]    <=  16'h783E;
                char10[13]    <=  16'h3FFE;
                char10[14]    <=  16'h0FDE;
                char10[15]    <=  16'h001C;
                char10[16]    <=  16'h003C;
                char10[17]    <=  16'h1838;
                char10[18]    <=  16'h3C78;
                char10[19]    <=  16'h3CF0;
                char10[20]    <=  16'h1FC0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end   
            default:begin
                char10[0]     <=  16'h0000;
                char10[1]     <=  16'h0000;
                char10[2]     <=  16'h0000;
                char10[3]     <=  16'h0000;
                char10[4]     <=  16'h07E0;
                char10[5]     <=  16'h0FF0;
                char10[6]     <=  16'h1C38;
                char10[7]     <=  16'h3C3C;
                char10[8]     <=  16'h781C;
                char10[9]     <=  16'h781E;
                char10[10]    <=  16'h781E;
                char10[11]    <=  16'h781E;
                char10[12]    <=  16'h781E;
                char10[13]    <=  16'h781E;
                char10[14]    <=  16'h781E;
                char10[15]    <=  16'h781E;
                char10[16]    <=  16'h781E;
                char10[17]    <=  16'h383C;
                char10[18]    <=  16'h3C38;
                char10[19]    <=  16'h1E78;
                char10[20]    <=  16'h07E0;
                char10[21]    <=  16'h0000;
                char10[22]    <=  16'h0000;
                char10[23]    <=  16'h0000;
            end
        endcase
always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char11[0]     <=  16'h0000;
       char11[1]     <=  16'h0000;
       char11[2]     <=  16'h0000;
       char11[3]     <=  16'h0000;
       char11[4]     <=  16'h07E0;
       char11[5]     <=  16'h0FF0;
       char11[6]     <=  16'h1C38;
       char11[7]     <=  16'h3C3C;
       char11[8]     <=  16'h781C;
       char11[9]     <=  16'h781E;
       char11[10]    <=  16'h781E;
       char11[11]    <=  16'h781E;
       char11[12]    <=  16'h781E;
       char11[13]    <=  16'h781E;
       char11[14]    <=  16'h781E;
       char11[15]    <=  16'h781E;
       char11[16]    <=  16'h781E;
       char11[17]    <=  16'h383C;
       char11[18]    <=  16'h3C38;
       char11[19]    <=  16'h1E78;
       char11[20]    <=  16'h07E0;
       char11[21]    <=  16'h0000;
       char11[22]    <=  16'h0000;
       char11[23]    <=  16'h0000;
    end
    else    
        case(ten2)
            4'd0  :  begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h07E0;
                char11[5]     <=  16'h0FF0;
                char11[6]     <=  16'h1C38;
                char11[7]     <=  16'h3C3C;
                char11[8]     <=  16'h781C;
                char11[9]     <=  16'h781E;
                char11[10]    <=  16'h781E;
                char11[11]    <=  16'h781E;
                char11[12]    <=  16'h781E;
                char11[13]    <=  16'h781E;
                char11[14]    <=  16'h781E;
                char11[15]    <=  16'h781E;
                char11[16]    <=  16'h781E;
                char11[17]    <=  16'h383C;
                char11[18]    <=  16'h3C38;
                char11[19]    <=  16'h1E78;
                char11[20]    <=  16'h07E0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h00C0;
                char11[5]     <=  16'h0FC0;
                char11[6]     <=  16'h1FC0;
                char11[7]     <=  16'h03C0;
                char11[8]     <=  16'h03C0;
                char11[9]     <=  16'h03C0;
                char11[10]    <=  16'h03C0;
                char11[11]    <=  16'h03C0;
                char11[12]    <=  16'h03C0;
                char11[13]    <=  16'h03C0;
                char11[14]    <=  16'h03C0;
                char11[15]    <=  16'h03C0;
                char11[16]    <=  16'h03C0;
                char11[17]    <=  16'h03C0;
                char11[18]    <=  16'h03C0;
                char11[19]    <=  16'h03E0;
                char11[20]    <=  16'h1FFC;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end
            4'd2  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h07E0;
                char11[5]     <=  16'h1EF8;
                char11[6]     <=  16'h383C;
                char11[7]     <=  16'h781C;
                char11[8]     <=  16'h7C1C;
                char11[9]     <=  16'h381C;
                char11[10]    <=  16'h003C;
                char11[11]    <=  16'h0038;
                char11[12]    <=  16'h0070;
                char11[13]    <=  16'h01E0;
                char11[14]    <=  16'h0380;
                char11[15]    <=  16'h0700;
                char11[16]    <=  16'h0E06;
                char11[17]    <=  16'h1C0E;
                char11[18]    <=  16'h301C;
                char11[19]    <=  16'h7FFC;
                char11[20]    <=  16'h7FFC;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h07E0;
                char11[5]     <=  16'h1EF0;
                char11[6]     <=  16'h3838;
                char11[7]     <=  16'h383C;
                char11[8]     <=  16'h383C;
                char11[9]     <=  16'h003C;
                char11[10]    <=  16'h0078;
                char11[11]    <=  16'h03F0;
                char11[12]    <=  16'h03F0;
                char11[13]    <=  16'h0038;
                char11[14]    <=  16'h001C;
                char11[15]    <=  16'h001E;
                char11[16]    <=  16'h381E;
                char11[17]    <=  16'h781E;
                char11[18]    <=  16'h783C;
                char11[19]    <=  16'h3C78;
                char11[20]    <=  16'h0FE0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h0070;
                char11[5]     <=  16'h0070;
                char11[6]     <=  16'h00F0;
                char11[7]     <=  16'h01F0;
                char11[8]     <=  16'h03F0;
                char11[9]     <=  16'h0770;
                char11[10]    <=  16'h0E70;
                char11[11]    <=  16'h0C70;
                char11[12]    <=  16'h1870;
                char11[13]    <=  16'h3070;
                char11[14]    <=  16'h7070;
                char11[15]    <=  16'hFFFF;
                char11[16]    <=  16'h0070;
                char11[17]    <=  16'h0070;
                char11[18]    <=  16'h0070;
                char11[19]    <=  16'h00F8;
                char11[20]    <=  16'h07FE;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h1FFC;
                char11[5]     <=  16'h1FFC;
                char11[6]     <=  16'h3800;
                char11[7]     <=  16'h3800;
                char11[8]     <=  16'h3800;
                char11[9]     <=  16'h3800;
                char11[10]    <=  16'h3FF0;
                char11[11]    <=  16'h3FF8;
                char11[12]    <=  16'h383C;
                char11[13]    <=  16'h101C;
                char11[14]    <=  16'h001E;
                char11[15]    <=  16'h001E;
                char11[16]    <=  16'h381E;
                char11[17]    <=  16'h781C;
                char11[18]    <=  16'h783C;
                char11[19]    <=  16'h3C78;
                char11[20]    <=  16'h0FF0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h03F0;
                char11[5]     <=  16'h0F38;
                char11[6]     <=  16'h1C3C;
                char11[7]     <=  16'h383C;
                char11[8]     <=  16'h3800;
                char11[9]     <=  16'h7800;
                char11[10]    <=  16'h7BF0;
                char11[11]    <=  16'h7FF8;
                char11[12]    <=  16'h7C3C;
                char11[13]    <=  16'h781E;
                char11[14]    <=  16'h781E;
                char11[15]    <=  16'h781E;
                char11[16]    <=  16'h781E;
                char11[17]    <=  16'h381E;
                char11[18]    <=  16'h3C1C;
                char11[19]    <=  16'h1E38;
                char11[20]    <=  16'h07F0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h3FFE;
                char11[5]     <=  16'h3FFE;
                char11[6]     <=  16'h381C;
                char11[7]     <=  16'h7018;
                char11[8]     <=  16'h7030;
                char11[9]     <=  16'h0070;
                char11[10]    <=  16'h00E0;
                char11[11]    <=  16'h00E0;
                char11[12]    <=  16'h01C0;
                char11[13]    <=  16'h01C0;
                char11[14]    <=  16'h0380;
                char11[15]    <=  16'h0380;
                char11[16]    <=  16'h0780;
                char11[17]    <=  16'h0780;
                char11[18]    <=  16'h0780;
                char11[19]    <=  16'h0780;
                char11[20]    <=  16'h0780;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h07E0;
                char11[5]     <=  16'h1E78;
                char11[6]     <=  16'h381C;
                char11[7]     <=  16'h701E;
                char11[8]     <=  16'h701E;
                char11[9]     <=  16'h781C;
                char11[10]    <=  16'h3E3C;
                char11[11]    <=  16'h1FF0;
                char11[12]    <=  16'h1FF0;
                char11[13]    <=  16'h3CF8;
                char11[14]    <=  16'h783C;
                char11[15]    <=  16'h701E;
                char11[16]    <=  16'h701E;
                char11[17]    <=  16'h701E;
                char11[18]    <=  16'h701C;
                char11[19]    <=  16'h3C38;
                char11[20]    <=  16'h0FF0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h0FE0;
                char11[5]     <=  16'h1EF8;
                char11[6]     <=  16'h3838;
                char11[7]     <=  16'h781C;
                char11[8]     <=  16'h701E;
                char11[9]     <=  16'h701E;
                char11[10]    <=  16'h701E;
                char11[11]    <=  16'h781E;
                char11[12]    <=  16'h783E;
                char11[13]    <=  16'h3FFE;
                char11[14]    <=  16'h0FDE;
                char11[15]    <=  16'h001C;
                char11[16]    <=  16'h003C;
                char11[17]    <=  16'h1838;
                char11[18]    <=  16'h3C78;
                char11[19]    <=  16'h3CF0;
                char11[20]    <=  16'h1FC0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end   
            default:begin
                char11[0]     <=  16'h0000;
                char11[1]     <=  16'h0000;
                char11[2]     <=  16'h0000;
                char11[3]     <=  16'h0000;
                char11[4]     <=  16'h07E0;
                char11[5]     <=  16'h0FF0;
                char11[6]     <=  16'h1C38;
                char11[7]     <=  16'h3C3C;
                char11[8]     <=  16'h781C;
                char11[9]     <=  16'h781E;
                char11[10]    <=  16'h781E;
                char11[11]    <=  16'h781E;
                char11[12]    <=  16'h781E;
                char11[13]    <=  16'h781E;
                char11[14]    <=  16'h781E;
                char11[15]    <=  16'h781E;
                char11[16]    <=  16'h781E;
                char11[17]    <=  16'h383C;
                char11[18]    <=  16'h3C38;
                char11[19]    <=  16'h1E78;
                char11[20]    <=  16'h07E0;
                char11[21]    <=  16'h0000;
                char11[22]    <=  16'h0000;
                char11[23]    <=  16'h0000;
            end
        endcase

always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char12[0]     <=  16'h0000;
       char12[1]     <=  16'h0000;
       char12[2]     <=  16'h0000;
       char12[3]     <=  16'h0000;
       char12[4]     <=  16'h07E0;
       char12[5]     <=  16'h0FF0;
       char12[6]     <=  16'h1C38;
       char12[7]     <=  16'h3C3C;
       char12[8]     <=  16'h781C;
       char12[9]     <=  16'h781E;
       char12[10]    <=  16'h781E;
       char12[11]    <=  16'h781E;
       char12[12]    <=  16'h781E;
       char12[13]    <=  16'h781E;
       char12[14]    <=  16'h781E;
       char12[15]    <=  16'h781E;
       char12[16]    <=  16'h781E;
       char12[17]    <=  16'h383C;
       char12[18]    <=  16'h3C38;
       char12[19]    <=  16'h1E78;
       char12[20]    <=  16'h07E0;
       char12[21]    <=  16'h0000;
       char12[22]    <=  16'h0000;
       char12[23]    <=  16'h0000;
    end
    else    
        case(unit2)
            4'd0  :  begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h07E0;
                char12[5]     <=  16'h0FF0;
                char12[6]     <=  16'h1C38;
                char12[7]     <=  16'h3C3C;
                char12[8]     <=  16'h781C;
                char12[9]     <=  16'h781E;
                char12[10]    <=  16'h781E;
                char12[11]    <=  16'h781E;
                char12[12]    <=  16'h781E;
                char12[13]    <=  16'h781E;
                char12[14]    <=  16'h781E;
                char12[15]    <=  16'h781E;
                char12[16]    <=  16'h781E;
                char12[17]    <=  16'h383C;
                char12[18]    <=  16'h3C38;
                char12[19]    <=  16'h1E78;
                char12[20]    <=  16'h07E0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h00C0;
                char12[5]     <=  16'h0FC0;
                char12[6]     <=  16'h1FC0;
                char12[7]     <=  16'h03C0;
                char12[8]     <=  16'h03C0;
                char12[9]     <=  16'h03C0;
                char12[10]    <=  16'h03C0;
                char12[11]    <=  16'h03C0;
                char12[12]    <=  16'h03C0;
                char12[13]    <=  16'h03C0;
                char12[14]    <=  16'h03C0;
                char12[15]    <=  16'h03C0;
                char12[16]    <=  16'h03C0;
                char12[17]    <=  16'h03C0;
                char12[18]    <=  16'h03C0;
                char12[19]    <=  16'h03E0;
                char12[20]    <=  16'h1FFC;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end
            4'd2  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h07E0;
                char12[5]     <=  16'h1EF8;
                char12[6]     <=  16'h383C;
                char12[7]     <=  16'h781C;
                char12[8]     <=  16'h7C1C;
                char12[9]     <=  16'h381C;
                char12[10]    <=  16'h003C;
                char12[11]    <=  16'h0038;
                char12[12]    <=  16'h0070;
                char12[13]    <=  16'h01E0;
                char12[14]    <=  16'h0380;
                char12[15]    <=  16'h0700;
                char12[16]    <=  16'h0E06;
                char12[17]    <=  16'h1C0E;
                char12[18]    <=  16'h301C;
                char12[19]    <=  16'h7FFC;
                char12[20]    <=  16'h7FFC;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h07E0;
                char12[5]     <=  16'h1EF0;
                char12[6]     <=  16'h3838;
                char12[7]     <=  16'h383C;
                char12[8]     <=  16'h383C;
                char12[9]     <=  16'h003C;
                char12[10]    <=  16'h0078;
                char12[11]    <=  16'h03F0;
                char12[12]    <=  16'h03F0;
                char12[13]    <=  16'h0038;
                char12[14]    <=  16'h001C;
                char12[15]    <=  16'h001E;
                char12[16]    <=  16'h381E;
                char12[17]    <=  16'h781E;
                char12[18]    <=  16'h783C;
                char12[19]    <=  16'h3C78;
                char12[20]    <=  16'h0FE0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h0070;
                char12[5]     <=  16'h0070;
                char12[6]     <=  16'h00F0;
                char12[7]     <=  16'h01F0;
                char12[8]     <=  16'h03F0;
                char12[9]     <=  16'h0770;
                char12[10]    <=  16'h0E70;
                char12[11]    <=  16'h0C70;
                char12[12]    <=  16'h1870;
                char12[13]    <=  16'h3070;
                char12[14]    <=  16'h7070;
                char12[15]    <=  16'hFFFF;
                char12[16]    <=  16'h0070;
                char12[17]    <=  16'h0070;
                char12[18]    <=  16'h0070;
                char12[19]    <=  16'h00F8;
                char12[20]    <=  16'h07FE;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h1FFC;
                char12[5]     <=  16'h1FFC;
                char12[6]     <=  16'h3800;
                char12[7]     <=  16'h3800;
                char12[8]     <=  16'h3800;
                char12[9]     <=  16'h3800;
                char12[10]    <=  16'h3FF0;
                char12[11]    <=  16'h3FF8;
                char12[12]    <=  16'h383C;
                char12[13]    <=  16'h101C;
                char12[14]    <=  16'h001E;
                char12[15]    <=  16'h001E;
                char12[16]    <=  16'h381E;
                char12[17]    <=  16'h781C;
                char12[18]    <=  16'h783C;
                char12[19]    <=  16'h3C78;
                char12[20]    <=  16'h0FF0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h03F0;
                char12[5]     <=  16'h0F38;
                char12[6]     <=  16'h1C3C;
                char12[7]     <=  16'h383C;
                char12[8]     <=  16'h3800;
                char12[9]     <=  16'h7800;
                char12[10]    <=  16'h7BF0;
                char12[11]    <=  16'h7FF8;
                char12[12]    <=  16'h7C3C;
                char12[13]    <=  16'h781E;
                char12[14]    <=  16'h781E;
                char12[15]    <=  16'h781E;
                char12[16]    <=  16'h781E;
                char12[17]    <=  16'h381E;
                char12[18]    <=  16'h3C1C;
                char12[19]    <=  16'h1E38;
                char12[20]    <=  16'h07F0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h3FFE;
                char12[5]     <=  16'h3FFE;
                char12[6]     <=  16'h381C;
                char12[7]     <=  16'h7018;
                char12[8]     <=  16'h7030;
                char12[9]     <=  16'h0070;
                char12[10]    <=  16'h00E0;
                char12[11]    <=  16'h00E0;
                char12[12]    <=  16'h01C0;
                char12[13]    <=  16'h01C0;
                char12[14]    <=  16'h0380;
                char12[15]    <=  16'h0380;
                char12[16]    <=  16'h0780;
                char12[17]    <=  16'h0780;
                char12[18]    <=  16'h0780;
                char12[19]    <=  16'h0780;
                char12[20]    <=  16'h0780;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h07E0;
                char12[5]     <=  16'h1E78;
                char12[6]     <=  16'h381C;
                char12[7]     <=  16'h701E;
                char12[8]     <=  16'h701E;
                char12[9]     <=  16'h781C;
                char12[10]    <=  16'h3E3C;
                char12[11]    <=  16'h1FF0;
                char12[12]    <=  16'h1FF0;
                char12[13]    <=  16'h3CF8;
                char12[14]    <=  16'h783C;
                char12[15]    <=  16'h701E;
                char12[16]    <=  16'h701E;
                char12[17]    <=  16'h701E;
                char12[18]    <=  16'h701C;
                char12[19]    <=  16'h3C38;
                char12[20]    <=  16'h0FF0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h0FE0;
                char12[5]     <=  16'h1EF8;
                char12[6]     <=  16'h3838;
                char12[7]     <=  16'h781C;
                char12[8]     <=  16'h701E;
                char12[9]     <=  16'h701E;
                char12[10]    <=  16'h701E;
                char12[11]    <=  16'h781E;
                char12[12]    <=  16'h783E;
                char12[13]    <=  16'h3FFE;
                char12[14]    <=  16'h0FDE;
                char12[15]    <=  16'h001C;
                char12[16]    <=  16'h003C;
                char12[17]    <=  16'h1838;
                char12[18]    <=  16'h3C78;
                char12[19]    <=  16'h3CF0;
                char12[20]    <=  16'h1FC0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end   
            default:begin
                char12[0]     <=  16'h0000;
                char12[1]     <=  16'h0000;
                char12[2]     <=  16'h0000;
                char12[3]     <=  16'h0000;
                char12[4]     <=  16'h07E0;
                char12[5]     <=  16'h0FF0;
                char12[6]     <=  16'h1C38;
                char12[7]     <=  16'h3C3C;
                char12[8]     <=  16'h781C;
                char12[9]     <=  16'h781E;
                char12[10]    <=  16'h781E;
                char12[11]    <=  16'h781E;
                char12[12]    <=  16'h781E;
                char12[13]    <=  16'h781E;
                char12[14]    <=  16'h781E;
                char12[15]    <=  16'h781E;
                char12[16]    <=  16'h781E;
                char12[17]    <=  16'h383C;
                char12[18]    <=  16'h3C38;
                char12[19]    <=  16'h1E78;
                char12[20]    <=  16'h07E0;
                char12[21]    <=  16'h0000;
                char12[22]    <=  16'h0000;
                char12[23]    <=  16'h0000;
            end
        endcase

//------------------------------------------------------------------------------
//--------------------------------------CH3-------------------------------------
//------------------------------------------------------------------------------



always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char13[0]     <=  16'h0000;
       char13[1]     <=  16'h0000;
       char13[2]     <=  16'h0000;
       char13[3]     <=  16'h0000;
       char13[4]     <=  16'h07E0;
       char13[5]     <=  16'h0FF0;
       char13[6]     <=  16'h1C38;
       char13[7]     <=  16'h3C3C;
       char13[8]     <=  16'h781C;
       char13[9]     <=  16'h781E;
       char13[10]    <=  16'h781E;
       char13[11]    <=  16'h781E;
       char13[12]    <=  16'h781E;
       char13[13]    <=  16'h781E;
       char13[14]    <=  16'h781E;
       char13[15]    <=  16'h781E;
       char13[16]    <=  16'h781E;
       char13[17]    <=  16'h383C;
       char13[18]    <=  16'h3C38;
       char13[19]    <=  16'h1E78;
       char13[20]    <=  16'h07E0;
       char13[21]    <=  16'h0000;
       char13[22]    <=  16'h0000;
       char13[23]    <=  16'h0000;
    end
    else    
        case(hun3)
            4'd0  :  begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h07E0;
                char13[5]     <=  16'h0FF0;
                char13[6]     <=  16'h1C38;
                char13[7]     <=  16'h3C3C;
                char13[8]     <=  16'h781C;
                char13[9]     <=  16'h781E;
                char13[10]    <=  16'h781E;
                char13[11]    <=  16'h781E;
                char13[12]    <=  16'h781E;
                char13[13]    <=  16'h781E;
                char13[14]    <=  16'h781E;
                char13[15]    <=  16'h781E;
                char13[16]    <=  16'h781E;
                char13[17]    <=  16'h383C;
                char13[18]    <=  16'h3C38;
                char13[19]    <=  16'h1E78;
                char13[20]    <=  16'h07E0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h00C0;
                char13[5]     <=  16'h0FC0;
                char13[6]     <=  16'h1FC0;
                char13[7]     <=  16'h03C0;
                char13[8]     <=  16'h03C0;
                char13[9]     <=  16'h03C0;
                char13[10]    <=  16'h03C0;
                char13[11]    <=  16'h03C0;
                char13[12]    <=  16'h03C0;
                char13[13]    <=  16'h03C0;
                char13[14]    <=  16'h03C0;
                char13[15]    <=  16'h03C0;
                char13[16]    <=  16'h03C0;
                char13[17]    <=  16'h03C0;
                char13[18]    <=  16'h03C0;
                char13[19]    <=  16'h03E0;
                char13[20]    <=  16'h1FFC;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end
            4'd2  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h07E0;
                char13[5]     <=  16'h1EF8;
                char13[6]     <=  16'h383C;
                char13[7]     <=  16'h781C;
                char13[8]     <=  16'h7C1C;
                char13[9]     <=  16'h381C;
                char13[10]    <=  16'h003C;
                char13[11]    <=  16'h0038;
                char13[12]    <=  16'h0070;
                char13[13]    <=  16'h01E0;
                char13[14]    <=  16'h0380;
                char13[15]    <=  16'h0700;
                char13[16]    <=  16'h0E06;
                char13[17]    <=  16'h1C0E;
                char13[18]    <=  16'h301C;
                char13[19]    <=  16'h7FFC;
                char13[20]    <=  16'h7FFC;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h07E0;
                char13[5]     <=  16'h1EF0;
                char13[6]     <=  16'h3838;
                char13[7]     <=  16'h383C;
                char13[8]     <=  16'h383C;
                char13[9]     <=  16'h003C;
                char13[10]    <=  16'h0078;
                char13[11]    <=  16'h03F0;
                char13[12]    <=  16'h03F0;
                char13[13]    <=  16'h0038;
                char13[14]    <=  16'h001C;
                char13[15]    <=  16'h001E;
                char13[16]    <=  16'h381E;
                char13[17]    <=  16'h781E;
                char13[18]    <=  16'h783C;
                char13[19]    <=  16'h3C78;
                char13[20]    <=  16'h0FE0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h0070;
                char13[5]     <=  16'h0070;
                char13[6]     <=  16'h00F0;
                char13[7]     <=  16'h01F0;
                char13[8]     <=  16'h03F0;
                char13[9]     <=  16'h0770;
                char13[10]    <=  16'h0E70;
                char13[11]    <=  16'h0C70;
                char13[12]    <=  16'h1870;
                char13[13]    <=  16'h3070;
                char13[14]    <=  16'h7070;
                char13[15]    <=  16'hFFFF;
                char13[16]    <=  16'h0070;
                char13[17]    <=  16'h0070;
                char13[18]    <=  16'h0070;
                char13[19]    <=  16'h00F8;
                char13[20]    <=  16'h07FE;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h1FFC;
                char13[5]     <=  16'h1FFC;
                char13[6]     <=  16'h3800;
                char13[7]     <=  16'h3800;
                char13[8]     <=  16'h3800;
                char13[9]     <=  16'h3800;
                char13[10]    <=  16'h3FF0;
                char13[11]    <=  16'h3FF8;
                char13[12]    <=  16'h383C;
                char13[13]    <=  16'h101C;
                char13[14]    <=  16'h001E;
                char13[15]    <=  16'h001E;
                char13[16]    <=  16'h381E;
                char13[17]    <=  16'h781C;
                char13[18]    <=  16'h783C;
                char13[19]    <=  16'h3C78;
                char13[20]    <=  16'h0FF0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h03F0;
                char13[5]     <=  16'h0F38;
                char13[6]     <=  16'h1C3C;
                char13[7]     <=  16'h383C;
                char13[8]     <=  16'h3800;
                char13[9]     <=  16'h7800;
                char13[10]    <=  16'h7BF0;
                char13[11]    <=  16'h7FF8;
                char13[12]    <=  16'h7C3C;
                char13[13]    <=  16'h781E;
                char13[14]    <=  16'h781E;
                char13[15]    <=  16'h781E;
                char13[16]    <=  16'h781E;
                char13[17]    <=  16'h381E;
                char13[18]    <=  16'h3C1C;
                char13[19]    <=  16'h1E38;
                char13[20]    <=  16'h07F0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h3FFE;
                char13[5]     <=  16'h3FFE;
                char13[6]     <=  16'h381C;
                char13[7]     <=  16'h7018;
                char13[8]     <=  16'h7030;
                char13[9]     <=  16'h0070;
                char13[10]    <=  16'h00E0;
                char13[11]    <=  16'h00E0;
                char13[12]    <=  16'h01C0;
                char13[13]    <=  16'h01C0;
                char13[14]    <=  16'h0380;
                char13[15]    <=  16'h0380;
                char13[16]    <=  16'h0780;
                char13[17]    <=  16'h0780;
                char13[18]    <=  16'h0780;
                char13[19]    <=  16'h0780;
                char13[20]    <=  16'h0780;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h07E0;
                char13[5]     <=  16'h1E78;
                char13[6]     <=  16'h381C;
                char13[7]     <=  16'h701E;
                char13[8]     <=  16'h701E;
                char13[9]     <=  16'h781C;
                char13[10]    <=  16'h3E3C;
                char13[11]    <=  16'h1FF0;
                char13[12]    <=  16'h1FF0;
                char13[13]    <=  16'h3CF8;
                char13[14]    <=  16'h783C;
                char13[15]    <=  16'h701E;
                char13[16]    <=  16'h701E;
                char13[17]    <=  16'h701E;
                char13[18]    <=  16'h701C;
                char13[19]    <=  16'h3C38;
                char13[20]    <=  16'h0FF0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h0FE0;
                char13[5]     <=  16'h1EF8;
                char13[6]     <=  16'h3838;
                char13[7]     <=  16'h781C;
                char13[8]     <=  16'h701E;
                char13[9]     <=  16'h701E;
                char13[10]    <=  16'h701E;
                char13[11]    <=  16'h781E;
                char13[12]    <=  16'h783E;
                char13[13]    <=  16'h3FFE;
                char13[14]    <=  16'h0FDE;
                char13[15]    <=  16'h001C;
                char13[16]    <=  16'h003C;
                char13[17]    <=  16'h1838;
                char13[18]    <=  16'h3C78;
                char13[19]    <=  16'h3CF0;
                char13[20]    <=  16'h1FC0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end   
            default:begin
                char13[0]     <=  16'h0000;
                char13[1]     <=  16'h0000;
                char13[2]     <=  16'h0000;
                char13[3]     <=  16'h0000;
                char13[4]     <=  16'h07E0;
                char13[5]     <=  16'h0FF0;
                char13[6]     <=  16'h1C38;
                char13[7]     <=  16'h3C3C;
                char13[8]     <=  16'h781C;
                char13[9]     <=  16'h781E;
                char13[10]    <=  16'h781E;
                char13[11]    <=  16'h781E;
                char13[12]    <=  16'h781E;
                char13[13]    <=  16'h781E;
                char13[14]    <=  16'h781E;
                char13[15]    <=  16'h781E;
                char13[16]    <=  16'h781E;
                char13[17]    <=  16'h383C;
                char13[18]    <=  16'h3C38;
                char13[19]    <=  16'h1E78;
                char13[20]    <=  16'h07E0;
                char13[21]    <=  16'h0000;
                char13[22]    <=  16'h0000;
                char13[23]    <=  16'h0000;
            end
        endcase
always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char14[0]     <=  16'h0000;
       char14[1]     <=  16'h0000;
       char14[2]     <=  16'h0000;
       char14[3]     <=  16'h0000;
       char14[4]     <=  16'h07E0;
       char14[5]     <=  16'h0FF0;
       char14[6]     <=  16'h1C38;
       char14[7]     <=  16'h3C3C;
       char14[8]     <=  16'h781C;
       char14[9]     <=  16'h781E;
       char14[10]    <=  16'h781E;
       char14[11]    <=  16'h781E;
       char14[12]    <=  16'h781E;
       char14[13]    <=  16'h781E;
       char14[14]    <=  16'h781E;
       char14[15]    <=  16'h781E;
       char14[16]    <=  16'h781E;
       char14[17]    <=  16'h383C;
       char14[18]    <=  16'h3C38;
       char14[19]    <=  16'h1E78;
       char14[20]    <=  16'h07E0;
       char14[21]    <=  16'h0000;
       char14[22]    <=  16'h0000;
       char14[23]    <=  16'h0000;
    end
    else    
        case(ten3)
            4'd0  :  begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h07E0;
                char14[5]     <=  16'h0FF0;
                char14[6]     <=  16'h1C38;
                char14[7]     <=  16'h3C3C;
                char14[8]     <=  16'h781C;
                char14[9]     <=  16'h781E;
                char14[10]    <=  16'h781E;
                char14[11]    <=  16'h781E;
                char14[12]    <=  16'h781E;
                char14[13]    <=  16'h781E;
                char14[14]    <=  16'h781E;
                char14[15]    <=  16'h781E;
                char14[16]    <=  16'h781E;
                char14[17]    <=  16'h383C;
                char14[18]    <=  16'h3C38;
                char14[19]    <=  16'h1E78;
                char14[20]    <=  16'h07E0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h00C0;
                char14[5]     <=  16'h0FC0;
                char14[6]     <=  16'h1FC0;
                char14[7]     <=  16'h03C0;
                char14[8]     <=  16'h03C0;
                char14[9]     <=  16'h03C0;
                char14[10]    <=  16'h03C0;
                char14[11]    <=  16'h03C0;
                char14[12]    <=  16'h03C0;
                char14[13]    <=  16'h03C0;
                char14[14]    <=  16'h03C0;
                char14[15]    <=  16'h03C0;
                char14[16]    <=  16'h03C0;
                char14[17]    <=  16'h03C0;
                char14[18]    <=  16'h03C0;
                char14[19]    <=  16'h03E0;
                char14[20]    <=  16'h1FFC;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end
            4'd2  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h07E0;
                char14[5]     <=  16'h1EF8;
                char14[6]     <=  16'h383C;
                char14[7]     <=  16'h781C;
                char14[8]     <=  16'h7C1C;
                char14[9]     <=  16'h381C;
                char14[10]    <=  16'h003C;
                char14[11]    <=  16'h0038;
                char14[12]    <=  16'h0070;
                char14[13]    <=  16'h01E0;
                char14[14]    <=  16'h0380;
                char14[15]    <=  16'h0700;
                char14[16]    <=  16'h0E06;
                char14[17]    <=  16'h1C0E;
                char14[18]    <=  16'h301C;
                char14[19]    <=  16'h7FFC;
                char14[20]    <=  16'h7FFC;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h07E0;
                char14[5]     <=  16'h1EF0;
                char14[6]     <=  16'h3838;
                char14[7]     <=  16'h383C;
                char14[8]     <=  16'h383C;
                char14[9]     <=  16'h003C;
                char14[10]    <=  16'h0078;
                char14[11]    <=  16'h03F0;
                char14[12]    <=  16'h03F0;
                char14[13]    <=  16'h0038;
                char14[14]    <=  16'h001C;
                char14[15]    <=  16'h001E;
                char14[16]    <=  16'h381E;
                char14[17]    <=  16'h781E;
                char14[18]    <=  16'h783C;
                char14[19]    <=  16'h3C78;
                char14[20]    <=  16'h0FE0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h0070;
                char14[5]     <=  16'h0070;
                char14[6]     <=  16'h00F0;
                char14[7]     <=  16'h01F0;
                char14[8]     <=  16'h03F0;
                char14[9]     <=  16'h0770;
                char14[10]    <=  16'h0E70;
                char14[11]    <=  16'h0C70;
                char14[12]    <=  16'h1870;
                char14[13]    <=  16'h3070;
                char14[14]    <=  16'h7070;
                char14[15]    <=  16'hFFFF;
                char14[16]    <=  16'h0070;
                char14[17]    <=  16'h0070;
                char14[18]    <=  16'h0070;
                char14[19]    <=  16'h00F8;
                char14[20]    <=  16'h07FE;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h1FFC;
                char14[5]     <=  16'h1FFC;
                char14[6]     <=  16'h3800;
                char14[7]     <=  16'h3800;
                char14[8]     <=  16'h3800;
                char14[9]     <=  16'h3800;
                char14[10]    <=  16'h3FF0;
                char14[11]    <=  16'h3FF8;
                char14[12]    <=  16'h383C;
                char14[13]    <=  16'h101C;
                char14[14]    <=  16'h001E;
                char14[15]    <=  16'h001E;
                char14[16]    <=  16'h381E;
                char14[17]    <=  16'h781C;
                char14[18]    <=  16'h783C;
                char14[19]    <=  16'h3C78;
                char14[20]    <=  16'h0FF0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h03F0;
                char14[5]     <=  16'h0F38;
                char14[6]     <=  16'h1C3C;
                char14[7]     <=  16'h383C;
                char14[8]     <=  16'h3800;
                char14[9]     <=  16'h7800;
                char14[10]    <=  16'h7BF0;
                char14[11]    <=  16'h7FF8;
                char14[12]    <=  16'h7C3C;
                char14[13]    <=  16'h781E;
                char14[14]    <=  16'h781E;
                char14[15]    <=  16'h781E;
                char14[16]    <=  16'h781E;
                char14[17]    <=  16'h381E;
                char14[18]    <=  16'h3C1C;
                char14[19]    <=  16'h1E38;
                char14[20]    <=  16'h07F0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h3FFE;
                char14[5]     <=  16'h3FFE;
                char14[6]     <=  16'h381C;
                char14[7]     <=  16'h7018;
                char14[8]     <=  16'h7030;
                char14[9]     <=  16'h0070;
                char14[10]    <=  16'h00E0;
                char14[11]    <=  16'h00E0;
                char14[12]    <=  16'h01C0;
                char14[13]    <=  16'h01C0;
                char14[14]    <=  16'h0380;
                char14[15]    <=  16'h0380;
                char14[16]    <=  16'h0780;
                char14[17]    <=  16'h0780;
                char14[18]    <=  16'h0780;
                char14[19]    <=  16'h0780;
                char14[20]    <=  16'h0780;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h07E0;
                char14[5]     <=  16'h1E78;
                char14[6]     <=  16'h381C;
                char14[7]     <=  16'h701E;
                char14[8]     <=  16'h701E;
                char14[9]     <=  16'h781C;
                char14[10]    <=  16'h3E3C;
                char14[11]    <=  16'h1FF0;
                char14[12]    <=  16'h1FF0;
                char14[13]    <=  16'h3CF8;
                char14[14]    <=  16'h783C;
                char14[15]    <=  16'h701E;
                char14[16]    <=  16'h701E;
                char14[17]    <=  16'h701E;
                char14[18]    <=  16'h701C;
                char14[19]    <=  16'h3C38;
                char14[20]    <=  16'h0FF0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h0FE0;
                char14[5]     <=  16'h1EF8;
                char14[6]     <=  16'h3838;
                char14[7]     <=  16'h781C;
                char14[8]     <=  16'h701E;
                char14[9]     <=  16'h701E;
                char14[10]    <=  16'h701E;
                char14[11]    <=  16'h781E;
                char14[12]    <=  16'h783E;
                char14[13]    <=  16'h3FFE;
                char14[14]    <=  16'h0FDE;
                char14[15]    <=  16'h001C;
                char14[16]    <=  16'h003C;
                char14[17]    <=  16'h1838;
                char14[18]    <=  16'h3C78;
                char14[19]    <=  16'h3CF0;
                char14[20]    <=  16'h1FC0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end   
            default:begin
                char14[0]     <=  16'h0000;
                char14[1]     <=  16'h0000;
                char14[2]     <=  16'h0000;
                char14[3]     <=  16'h0000;
                char14[4]     <=  16'h07E0;
                char14[5]     <=  16'h0FF0;
                char14[6]     <=  16'h1C38;
                char14[7]     <=  16'h3C3C;
                char14[8]     <=  16'h781C;
                char14[9]     <=  16'h781E;
                char14[10]    <=  16'h781E;
                char14[11]    <=  16'h781E;
                char14[12]    <=  16'h781E;
                char14[13]    <=  16'h781E;
                char14[14]    <=  16'h781E;
                char14[15]    <=  16'h781E;
                char14[16]    <=  16'h781E;
                char14[17]    <=  16'h383C;
                char14[18]    <=  16'h3C38;
                char14[19]    <=  16'h1E78;
                char14[20]    <=  16'h07E0;
                char14[21]    <=  16'h0000;
                char14[22]    <=  16'h0000;
                char14[23]    <=  16'h0000;
            end
        endcase

always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char15[0]     <=  16'h0000;
       char15[1]     <=  16'h0000;
       char15[2]     <=  16'h0000;
       char15[3]     <=  16'h0000;
       char15[4]     <=  16'h07E0;
       char15[5]     <=  16'h0FF0;
       char15[6]     <=  16'h1C38;
       char15[7]     <=  16'h3C3C;
       char15[8]     <=  16'h781C;
       char15[9]     <=  16'h781E;
       char15[10]    <=  16'h781E;
       char15[11]    <=  16'h781E;
       char15[12]    <=  16'h781E;
       char15[13]    <=  16'h781E;
       char15[14]    <=  16'h781E;
       char15[15]    <=  16'h781E;
       char15[16]    <=  16'h781E;
       char15[17]    <=  16'h383C;
       char15[18]    <=  16'h3C38;
       char15[19]    <=  16'h1E78;
       char15[20]    <=  16'h07E0;
       char15[21]    <=  16'h0000;
       char15[22]    <=  16'h0000;
       char15[23]    <=  16'h0000;
    end
    else    
        case(unit3)
            4'd0  :  begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h07E0;
                char15[5]     <=  16'h0FF0;
                char15[6]     <=  16'h1C38;
                char15[7]     <=  16'h3C3C;
                char15[8]     <=  16'h781C;
                char15[9]     <=  16'h781E;
                char15[10]    <=  16'h781E;
                char15[11]    <=  16'h781E;
                char15[12]    <=  16'h781E;
                char15[13]    <=  16'h781E;
                char15[14]    <=  16'h781E;
                char15[15]    <=  16'h781E;
                char15[16]    <=  16'h781E;
                char15[17]    <=  16'h383C;
                char15[18]    <=  16'h3C38;
                char15[19]    <=  16'h1E78;
                char15[20]    <=  16'h07E0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h00C0;
                char15[5]     <=  16'h0FC0;
                char15[6]     <=  16'h1FC0;
                char15[7]     <=  16'h03C0;
                char15[8]     <=  16'h03C0;
                char15[9]     <=  16'h03C0;
                char15[10]    <=  16'h03C0;
                char15[11]    <=  16'h03C0;
                char15[12]    <=  16'h03C0;
                char15[13]    <=  16'h03C0;
                char15[14]    <=  16'h03C0;
                char15[15]    <=  16'h03C0;
                char15[16]    <=  16'h03C0;
                char15[17]    <=  16'h03C0;
                char15[18]    <=  16'h03C0;
                char15[19]    <=  16'h03E0;
                char15[20]    <=  16'h1FFC;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end
            4'd2  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h07E0;
                char15[5]     <=  16'h1EF8;
                char15[6]     <=  16'h383C;
                char15[7]     <=  16'h781C;
                char15[8]     <=  16'h7C1C;
                char15[9]     <=  16'h381C;
                char15[10]    <=  16'h003C;
                char15[11]    <=  16'h0038;
                char15[12]    <=  16'h0070;
                char15[13]    <=  16'h01E0;
                char15[14]    <=  16'h0380;
                char15[15]    <=  16'h0700;
                char15[16]    <=  16'h0E06;
                char15[17]    <=  16'h1C0E;
                char15[18]    <=  16'h301C;
                char15[19]    <=  16'h7FFC;
                char15[20]    <=  16'h7FFC;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h07E0;
                char15[5]     <=  16'h1EF0;
                char15[6]     <=  16'h3838;
                char15[7]     <=  16'h383C;
                char15[8]     <=  16'h383C;
                char15[9]     <=  16'h003C;
                char15[10]    <=  16'h0078;
                char15[11]    <=  16'h03F0;
                char15[12]    <=  16'h03F0;
                char15[13]    <=  16'h0038;
                char15[14]    <=  16'h001C;
                char15[15]    <=  16'h001E;
                char15[16]    <=  16'h381E;
                char15[17]    <=  16'h781E;
                char15[18]    <=  16'h783C;
                char15[19]    <=  16'h3C78;
                char15[20]    <=  16'h0FE0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h0070;
                char15[5]     <=  16'h0070;
                char15[6]     <=  16'h00F0;
                char15[7]     <=  16'h01F0;
                char15[8]     <=  16'h03F0;
                char15[9]     <=  16'h0770;
                char15[10]    <=  16'h0E70;
                char15[11]    <=  16'h0C70;
                char15[12]    <=  16'h1870;
                char15[13]    <=  16'h3070;
                char15[14]    <=  16'h7070;
                char15[15]    <=  16'hFFFF;
                char15[16]    <=  16'h0070;
                char15[17]    <=  16'h0070;
                char15[18]    <=  16'h0070;
                char15[19]    <=  16'h00F8;
                char15[20]    <=  16'h07FE;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h1FFC;
                char15[5]     <=  16'h1FFC;
                char15[6]     <=  16'h3800;
                char15[7]     <=  16'h3800;
                char15[8]     <=  16'h3800;
                char15[9]     <=  16'h3800;
                char15[10]    <=  16'h3FF0;
                char15[11]    <=  16'h3FF8;
                char15[12]    <=  16'h383C;
                char15[13]    <=  16'h101C;
                char15[14]    <=  16'h001E;
                char15[15]    <=  16'h001E;
                char15[16]    <=  16'h381E;
                char15[17]    <=  16'h781C;
                char15[18]    <=  16'h783C;
                char15[19]    <=  16'h3C78;
                char15[20]    <=  16'h0FF0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h03F0;
                char15[5]     <=  16'h0F38;
                char15[6]     <=  16'h1C3C;
                char15[7]     <=  16'h383C;
                char15[8]     <=  16'h3800;
                char15[9]     <=  16'h7800;
                char15[10]    <=  16'h7BF0;
                char15[11]    <=  16'h7FF8;
                char15[12]    <=  16'h7C3C;
                char15[13]    <=  16'h781E;
                char15[14]    <=  16'h781E;
                char15[15]    <=  16'h781E;
                char15[16]    <=  16'h781E;
                char15[17]    <=  16'h381E;
                char15[18]    <=  16'h3C1C;
                char15[19]    <=  16'h1E38;
                char15[20]    <=  16'h07F0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h3FFE;
                char15[5]     <=  16'h3FFE;
                char15[6]     <=  16'h381C;
                char15[7]     <=  16'h7018;
                char15[8]     <=  16'h7030;
                char15[9]     <=  16'h0070;
                char15[10]    <=  16'h00E0;
                char15[11]    <=  16'h00E0;
                char15[12]    <=  16'h01C0;
                char15[13]    <=  16'h01C0;
                char15[14]    <=  16'h0380;
                char15[15]    <=  16'h0380;
                char15[16]    <=  16'h0780;
                char15[17]    <=  16'h0780;
                char15[18]    <=  16'h0780;
                char15[19]    <=  16'h0780;
                char15[20]    <=  16'h0780;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h07E0;
                char15[5]     <=  16'h1E78;
                char15[6]     <=  16'h381C;
                char15[7]     <=  16'h701E;
                char15[8]     <=  16'h701E;
                char15[9]     <=  16'h781C;
                char15[10]    <=  16'h3E3C;
                char15[11]    <=  16'h1FF0;
                char15[12]    <=  16'h1FF0;
                char15[13]    <=  16'h3CF8;
                char15[14]    <=  16'h783C;
                char15[15]    <=  16'h701E;
                char15[16]    <=  16'h701E;
                char15[17]    <=  16'h701E;
                char15[18]    <=  16'h701C;
                char15[19]    <=  16'h3C38;
                char15[20]    <=  16'h0FF0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h0FE0;
                char15[5]     <=  16'h1EF8;
                char15[6]     <=  16'h3838;
                char15[7]     <=  16'h781C;
                char15[8]     <=  16'h701E;
                char15[9]     <=  16'h701E;
                char15[10]    <=  16'h701E;
                char15[11]    <=  16'h781E;
                char15[12]    <=  16'h783E;
                char15[13]    <=  16'h3FFE;
                char15[14]    <=  16'h0FDE;
                char15[15]    <=  16'h001C;
                char15[16]    <=  16'h003C;
                char15[17]    <=  16'h1838;
                char15[18]    <=  16'h3C78;
                char15[19]    <=  16'h3CF0;
                char15[20]    <=  16'h1FC0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end   
            default:begin
                char15[0]     <=  16'h0000;
                char15[1]     <=  16'h0000;
                char15[2]     <=  16'h0000;
                char15[3]     <=  16'h0000;
                char15[4]     <=  16'h07E0;
                char15[5]     <=  16'h0FF0;
                char15[6]     <=  16'h1C38;
                char15[7]     <=  16'h3C3C;
                char15[8]     <=  16'h781C;
                char15[9]     <=  16'h781E;
                char15[10]    <=  16'h781E;
                char15[11]    <=  16'h781E;
                char15[12]    <=  16'h781E;
                char15[13]    <=  16'h781E;
                char15[14]    <=  16'h781E;
                char15[15]    <=  16'h781E;
                char15[16]    <=  16'h781E;
                char15[17]    <=  16'h383C;
                char15[18]    <=  16'h3C38;
                char15[19]    <=  16'h1E78;
                char15[20]    <=  16'h07E0;
                char15[21]    <=  16'h0000;
                char15[22]    <=  16'h0000;
                char15[23]    <=  16'h0000;
            end
        endcase

//------------------------------------------------------------------------------
//--------------------------------------CH4-------------------------------------
//------------------------------------------------------------------------------



always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char16[0]     <=  16'h0000;
       char16[1]     <=  16'h0000;
       char16[2]     <=  16'h0000;
       char16[3]     <=  16'h0000;
       char16[4]     <=  16'h07E0;
       char16[5]     <=  16'h0FF0;
       char16[6]     <=  16'h1C38;
       char16[7]     <=  16'h3C3C;
       char16[8]     <=  16'h781C;
       char16[9]     <=  16'h781E;
       char16[10]    <=  16'h781E;
       char16[11]    <=  16'h781E;
       char16[12]    <=  16'h781E;
       char16[13]    <=  16'h781E;
       char16[14]    <=  16'h781E;
       char16[15]    <=  16'h781E;
       char16[16]    <=  16'h781E;
       char16[17]    <=  16'h383C;
       char16[18]    <=  16'h3C38;
       char16[19]    <=  16'h1E78;
       char16[20]    <=  16'h07E0;
       char16[21]    <=  16'h0000;
       char16[22]    <=  16'h0000;
       char16[23]    <=  16'h0000;
    end
    else    
        case(hun4)
            4'd0  :  begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h07E0;
                char16[5]     <=  16'h0FF0;
                char16[6]     <=  16'h1C38;
                char16[7]     <=  16'h3C3C;
                char16[8]     <=  16'h781C;
                char16[9]     <=  16'h781E;
                char16[10]    <=  16'h781E;
                char16[11]    <=  16'h781E;
                char16[12]    <=  16'h781E;
                char16[13]    <=  16'h781E;
                char16[14]    <=  16'h781E;
                char16[15]    <=  16'h781E;
                char16[16]    <=  16'h781E;
                char16[17]    <=  16'h383C;
                char16[18]    <=  16'h3C38;
                char16[19]    <=  16'h1E78;
                char16[20]    <=  16'h07E0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h00C0;
                char16[5]     <=  16'h0FC0;
                char16[6]     <=  16'h1FC0;
                char16[7]     <=  16'h03C0;
                char16[8]     <=  16'h03C0;
                char16[9]     <=  16'h03C0;
                char16[10]    <=  16'h03C0;
                char16[11]    <=  16'h03C0;
                char16[12]    <=  16'h03C0;
                char16[13]    <=  16'h03C0;
                char16[14]    <=  16'h03C0;
                char16[15]    <=  16'h03C0;
                char16[16]    <=  16'h03C0;
                char16[17]    <=  16'h03C0;
                char16[18]    <=  16'h03C0;
                char16[19]    <=  16'h03E0;
                char16[20]    <=  16'h1FFC;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end
            4'd2  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h07E0;
                char16[5]     <=  16'h1EF8;
                char16[6]     <=  16'h383C;
                char16[7]     <=  16'h781C;
                char16[8]     <=  16'h7C1C;
                char16[9]     <=  16'h381C;
                char16[10]    <=  16'h003C;
                char16[11]    <=  16'h0038;
                char16[12]    <=  16'h0070;
                char16[13]    <=  16'h01E0;
                char16[14]    <=  16'h0380;
                char16[15]    <=  16'h0700;
                char16[16]    <=  16'h0E06;
                char16[17]    <=  16'h1C0E;
                char16[18]    <=  16'h301C;
                char16[19]    <=  16'h7FFC;
                char16[20]    <=  16'h7FFC;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h07E0;
                char16[5]     <=  16'h1EF0;
                char16[6]     <=  16'h3838;
                char16[7]     <=  16'h383C;
                char16[8]     <=  16'h383C;
                char16[9]     <=  16'h003C;
                char16[10]    <=  16'h0078;
                char16[11]    <=  16'h03F0;
                char16[12]    <=  16'h03F0;
                char16[13]    <=  16'h0038;
                char16[14]    <=  16'h001C;
                char16[15]    <=  16'h001E;
                char16[16]    <=  16'h381E;
                char16[17]    <=  16'h781E;
                char16[18]    <=  16'h783C;
                char16[19]    <=  16'h3C78;
                char16[20]    <=  16'h0FE0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h0070;
                char16[5]     <=  16'h0070;
                char16[6]     <=  16'h00F0;
                char16[7]     <=  16'h01F0;
                char16[8]     <=  16'h03F0;
                char16[9]     <=  16'h0770;
                char16[10]    <=  16'h0E70;
                char16[11]    <=  16'h0C70;
                char16[12]    <=  16'h1870;
                char16[13]    <=  16'h3070;
                char16[14]    <=  16'h7070;
                char16[15]    <=  16'hFFFF;
                char16[16]    <=  16'h0070;
                char16[17]    <=  16'h0070;
                char16[18]    <=  16'h0070;
                char16[19]    <=  16'h00F8;
                char16[20]    <=  16'h07FE;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h1FFC;
                char16[5]     <=  16'h1FFC;
                char16[6]     <=  16'h3800;
                char16[7]     <=  16'h3800;
                char16[8]     <=  16'h3800;
                char16[9]     <=  16'h3800;
                char16[10]    <=  16'h3FF0;
                char16[11]    <=  16'h3FF8;
                char16[12]    <=  16'h383C;
                char16[13]    <=  16'h101C;
                char16[14]    <=  16'h001E;
                char16[15]    <=  16'h001E;
                char16[16]    <=  16'h381E;
                char16[17]    <=  16'h781C;
                char16[18]    <=  16'h783C;
                char16[19]    <=  16'h3C78;
                char16[20]    <=  16'h0FF0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h03F0;
                char16[5]     <=  16'h0F38;
                char16[6]     <=  16'h1C3C;
                char16[7]     <=  16'h383C;
                char16[8]     <=  16'h3800;
                char16[9]     <=  16'h7800;
                char16[10]    <=  16'h7BF0;
                char16[11]    <=  16'h7FF8;
                char16[12]    <=  16'h7C3C;
                char16[13]    <=  16'h781E;
                char16[14]    <=  16'h781E;
                char16[15]    <=  16'h781E;
                char16[16]    <=  16'h781E;
                char16[17]    <=  16'h381E;
                char16[18]    <=  16'h3C1C;
                char16[19]    <=  16'h1E38;
                char16[20]    <=  16'h07F0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h3FFE;
                char16[5]     <=  16'h3FFE;
                char16[6]     <=  16'h381C;
                char16[7]     <=  16'h7018;
                char16[8]     <=  16'h7030;
                char16[9]     <=  16'h0070;
                char16[10]    <=  16'h00E0;
                char16[11]    <=  16'h00E0;
                char16[12]    <=  16'h01C0;
                char16[13]    <=  16'h01C0;
                char16[14]    <=  16'h0380;
                char16[15]    <=  16'h0380;
                char16[16]    <=  16'h0780;
                char16[17]    <=  16'h0780;
                char16[18]    <=  16'h0780;
                char16[19]    <=  16'h0780;
                char16[20]    <=  16'h0780;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h07E0;
                char16[5]     <=  16'h1E78;
                char16[6]     <=  16'h381C;
                char16[7]     <=  16'h701E;
                char16[8]     <=  16'h701E;
                char16[9]     <=  16'h781C;
                char16[10]    <=  16'h3E3C;
                char16[11]    <=  16'h1FF0;
                char16[12]    <=  16'h1FF0;
                char16[13]    <=  16'h3CF8;
                char16[14]    <=  16'h783C;
                char16[15]    <=  16'h701E;
                char16[16]    <=  16'h701E;
                char16[17]    <=  16'h701E;
                char16[18]    <=  16'h701C;
                char16[19]    <=  16'h3C38;
                char16[20]    <=  16'h0FF0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h0FE0;
                char16[5]     <=  16'h1EF8;
                char16[6]     <=  16'h3838;
                char16[7]     <=  16'h781C;
                char16[8]     <=  16'h701E;
                char16[9]     <=  16'h701E;
                char16[10]    <=  16'h701E;
                char16[11]    <=  16'h781E;
                char16[12]    <=  16'h783E;
                char16[13]    <=  16'h3FFE;
                char16[14]    <=  16'h0FDE;
                char16[15]    <=  16'h001C;
                char16[16]    <=  16'h003C;
                char16[17]    <=  16'h1838;
                char16[18]    <=  16'h3C78;
                char16[19]    <=  16'h3CF0;
                char16[20]    <=  16'h1FC0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end   
            default:begin
                char16[0]     <=  16'h0000;
                char16[1]     <=  16'h0000;
                char16[2]     <=  16'h0000;
                char16[3]     <=  16'h0000;
                char16[4]     <=  16'h07E0;
                char16[5]     <=  16'h0FF0;
                char16[6]     <=  16'h1C38;
                char16[7]     <=  16'h3C3C;
                char16[8]     <=  16'h781C;
                char16[9]     <=  16'h781E;
                char16[10]    <=  16'h781E;
                char16[11]    <=  16'h781E;
                char16[12]    <=  16'h781E;
                char16[13]    <=  16'h781E;
                char16[14]    <=  16'h781E;
                char16[15]    <=  16'h781E;
                char16[16]    <=  16'h781E;
                char16[17]    <=  16'h383C;
                char16[18]    <=  16'h3C38;
                char16[19]    <=  16'h1E78;
                char16[20]    <=  16'h07E0;
                char16[21]    <=  16'h0000;
                char16[22]    <=  16'h0000;
                char16[23]    <=  16'h0000;
            end
        endcase
always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char17[0]     <=  16'h0000;
       char17[1]     <=  16'h0000;
       char17[2]     <=  16'h0000;
       char17[3]     <=  16'h0000;
       char17[4]     <=  16'h07E0;
       char17[5]     <=  16'h0FF0;
       char17[6]     <=  16'h1C38;
       char17[7]     <=  16'h3C3C;
       char17[8]     <=  16'h781C;
       char17[9]     <=  16'h781E;
       char17[10]    <=  16'h781E;
       char17[11]    <=  16'h781E;
       char17[12]    <=  16'h781E;
       char17[13]    <=  16'h781E;
       char17[14]    <=  16'h781E;
       char17[15]    <=  16'h781E;
       char17[16]    <=  16'h781E;
       char17[17]    <=  16'h383C;
       char17[18]    <=  16'h3C38;
       char17[19]    <=  16'h1E78;
       char17[20]    <=  16'h07E0;
       char17[21]    <=  16'h0000;
       char17[22]    <=  16'h0000;
       char17[23]    <=  16'h0000;
    end
    else    
        case(ten4)
            4'd0  :  begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h07E0;
                char17[5]     <=  16'h0FF0;
                char17[6]     <=  16'h1C38;
                char17[7]     <=  16'h3C3C;
                char17[8]     <=  16'h781C;
                char17[9]     <=  16'h781E;
                char17[10]    <=  16'h781E;
                char17[11]    <=  16'h781E;
                char17[12]    <=  16'h781E;
                char17[13]    <=  16'h781E;
                char17[14]    <=  16'h781E;
                char17[15]    <=  16'h781E;
                char17[16]    <=  16'h781E;
                char17[17]    <=  16'h383C;
                char17[18]    <=  16'h3C38;
                char17[19]    <=  16'h1E78;
                char17[20]    <=  16'h07E0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h00C0;
                char17[5]     <=  16'h0FC0;
                char17[6]     <=  16'h1FC0;
                char17[7]     <=  16'h03C0;
                char17[8]     <=  16'h03C0;
                char17[9]     <=  16'h03C0;
                char17[10]    <=  16'h03C0;
                char17[11]    <=  16'h03C0;
                char17[12]    <=  16'h03C0;
                char17[13]    <=  16'h03C0;
                char17[14]    <=  16'h03C0;
                char17[15]    <=  16'h03C0;
                char17[16]    <=  16'h03C0;
                char17[17]    <=  16'h03C0;
                char17[18]    <=  16'h03C0;
                char17[19]    <=  16'h03E0;
                char17[20]    <=  16'h1FFC;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end
            4'd2  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h07E0;
                char17[5]     <=  16'h1EF8;
                char17[6]     <=  16'h383C;
                char17[7]     <=  16'h781C;
                char17[8]     <=  16'h7C1C;
                char17[9]     <=  16'h381C;
                char17[10]    <=  16'h003C;
                char17[11]    <=  16'h0038;
                char17[12]    <=  16'h0070;
                char17[13]    <=  16'h01E0;
                char17[14]    <=  16'h0380;
                char17[15]    <=  16'h0700;
                char17[16]    <=  16'h0E06;
                char17[17]    <=  16'h1C0E;
                char17[18]    <=  16'h301C;
                char17[19]    <=  16'h7FFC;
                char17[20]    <=  16'h7FFC;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h07E0;
                char17[5]     <=  16'h1EF0;
                char17[6]     <=  16'h3838;
                char17[7]     <=  16'h383C;
                char17[8]     <=  16'h383C;
                char17[9]     <=  16'h003C;
                char17[10]    <=  16'h0078;
                char17[11]    <=  16'h03F0;
                char17[12]    <=  16'h03F0;
                char17[13]    <=  16'h0038;
                char17[14]    <=  16'h001C;
                char17[15]    <=  16'h001E;
                char17[16]    <=  16'h381E;
                char17[17]    <=  16'h781E;
                char17[18]    <=  16'h783C;
                char17[19]    <=  16'h3C78;
                char17[20]    <=  16'h0FE0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h0070;
                char17[5]     <=  16'h0070;
                char17[6]     <=  16'h00F0;
                char17[7]     <=  16'h01F0;
                char17[8]     <=  16'h03F0;
                char17[9]     <=  16'h0770;
                char17[10]    <=  16'h0E70;
                char17[11]    <=  16'h0C70;
                char17[12]    <=  16'h1870;
                char17[13]    <=  16'h3070;
                char17[14]    <=  16'h7070;
                char17[15]    <=  16'hFFFF;
                char17[16]    <=  16'h0070;
                char17[17]    <=  16'h0070;
                char17[18]    <=  16'h0070;
                char17[19]    <=  16'h00F8;
                char17[20]    <=  16'h07FE;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h1FFC;
                char17[5]     <=  16'h1FFC;
                char17[6]     <=  16'h3800;
                char17[7]     <=  16'h3800;
                char17[8]     <=  16'h3800;
                char17[9]     <=  16'h3800;
                char17[10]    <=  16'h3FF0;
                char17[11]    <=  16'h3FF8;
                char17[12]    <=  16'h383C;
                char17[13]    <=  16'h101C;
                char17[14]    <=  16'h001E;
                char17[15]    <=  16'h001E;
                char17[16]    <=  16'h381E;
                char17[17]    <=  16'h781C;
                char17[18]    <=  16'h783C;
                char17[19]    <=  16'h3C78;
                char17[20]    <=  16'h0FF0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h03F0;
                char17[5]     <=  16'h0F38;
                char17[6]     <=  16'h1C3C;
                char17[7]     <=  16'h383C;
                char17[8]     <=  16'h3800;
                char17[9]     <=  16'h7800;
                char17[10]    <=  16'h7BF0;
                char17[11]    <=  16'h7FF8;
                char17[12]    <=  16'h7C3C;
                char17[13]    <=  16'h781E;
                char17[14]    <=  16'h781E;
                char17[15]    <=  16'h781E;
                char17[16]    <=  16'h781E;
                char17[17]    <=  16'h381E;
                char17[18]    <=  16'h3C1C;
                char17[19]    <=  16'h1E38;
                char17[20]    <=  16'h07F0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h3FFE;
                char17[5]     <=  16'h3FFE;
                char17[6]     <=  16'h381C;
                char17[7]     <=  16'h7018;
                char17[8]     <=  16'h7030;
                char17[9]     <=  16'h0070;
                char17[10]    <=  16'h00E0;
                char17[11]    <=  16'h00E0;
                char17[12]    <=  16'h01C0;
                char17[13]    <=  16'h01C0;
                char17[14]    <=  16'h0380;
                char17[15]    <=  16'h0380;
                char17[16]    <=  16'h0780;
                char17[17]    <=  16'h0780;
                char17[18]    <=  16'h0780;
                char17[19]    <=  16'h0780;
                char17[20]    <=  16'h0780;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h07E0;
                char17[5]     <=  16'h1E78;
                char17[6]     <=  16'h381C;
                char17[7]     <=  16'h701E;
                char17[8]     <=  16'h701E;
                char17[9]     <=  16'h781C;
                char17[10]    <=  16'h3E3C;
                char17[11]    <=  16'h1FF0;
                char17[12]    <=  16'h1FF0;
                char17[13]    <=  16'h3CF8;
                char17[14]    <=  16'h783C;
                char17[15]    <=  16'h701E;
                char17[16]    <=  16'h701E;
                char17[17]    <=  16'h701E;
                char17[18]    <=  16'h701C;
                char17[19]    <=  16'h3C38;
                char17[20]    <=  16'h0FF0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h0FE0;
                char17[5]     <=  16'h1EF8;
                char17[6]     <=  16'h3838;
                char17[7]     <=  16'h781C;
                char17[8]     <=  16'h701E;
                char17[9]     <=  16'h701E;
                char17[10]    <=  16'h701E;
                char17[11]    <=  16'h781E;
                char17[12]    <=  16'h783E;
                char17[13]    <=  16'h3FFE;
                char17[14]    <=  16'h0FDE;
                char17[15]    <=  16'h001C;
                char17[16]    <=  16'h003C;
                char17[17]    <=  16'h1838;
                char17[18]    <=  16'h3C78;
                char17[19]    <=  16'h3CF0;
                char17[20]    <=  16'h1FC0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end   
            default:begin
                char17[0]     <=  16'h0000;
                char17[1]     <=  16'h0000;
                char17[2]     <=  16'h0000;
                char17[3]     <=  16'h0000;
                char17[4]     <=  16'h07E0;
                char17[5]     <=  16'h0FF0;
                char17[6]     <=  16'h1C38;
                char17[7]     <=  16'h3C3C;
                char17[8]     <=  16'h781C;
                char17[9]     <=  16'h781E;
                char17[10]    <=  16'h781E;
                char17[11]    <=  16'h781E;
                char17[12]    <=  16'h781E;
                char17[13]    <=  16'h781E;
                char17[14]    <=  16'h781E;
                char17[15]    <=  16'h781E;
                char17[16]    <=  16'h781E;
                char17[17]    <=  16'h383C;
                char17[18]    <=  16'h3C38;
                char17[19]    <=  16'h1E78;
                char17[20]    <=  16'h07E0;
                char17[21]    <=  16'h0000;
                char17[22]    <=  16'h0000;
                char17[23]    <=  16'h0000;
            end
        endcase

always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char18[0]     <=  16'h0000;
       char18[1]     <=  16'h0000;
       char18[2]     <=  16'h0000;
       char18[3]     <=  16'h0000;
       char18[4]     <=  16'h07E0;
       char18[5]     <=  16'h0FF0;
       char18[6]     <=  16'h1C38;
       char18[7]     <=  16'h3C3C;
       char18[8]     <=  16'h781C;
       char18[9]     <=  16'h781E;
       char18[10]    <=  16'h781E;
       char18[11]    <=  16'h781E;
       char18[12]    <=  16'h781E;
       char18[13]    <=  16'h781E;
       char18[14]    <=  16'h781E;
       char18[15]    <=  16'h781E;
       char18[16]    <=  16'h781E;
       char18[17]    <=  16'h383C;
       char18[18]    <=  16'h3C38;
       char18[19]    <=  16'h1E78;
       char18[20]    <=  16'h07E0;
       char18[21]    <=  16'h0000;
       char18[22]    <=  16'h0000;
       char18[23]    <=  16'h0000;
    end
    else    
        case(unit4)
            4'd0  :  begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h07E0;
                char18[5]     <=  16'h0FF0;
                char18[6]     <=  16'h1C38;
                char18[7]     <=  16'h3C3C;
                char18[8]     <=  16'h781C;
                char18[9]     <=  16'h781E;
                char18[10]    <=  16'h781E;
                char18[11]    <=  16'h781E;
                char18[12]    <=  16'h781E;
                char18[13]    <=  16'h781E;
                char18[14]    <=  16'h781E;
                char18[15]    <=  16'h781E;
                char18[16]    <=  16'h781E;
                char18[17]    <=  16'h383C;
                char18[18]    <=  16'h3C38;
                char18[19]    <=  16'h1E78;
                char18[20]    <=  16'h07E0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h00C0;
                char18[5]     <=  16'h0FC0;
                char18[6]     <=  16'h1FC0;
                char18[7]     <=  16'h03C0;
                char18[8]     <=  16'h03C0;
                char18[9]     <=  16'h03C0;
                char18[10]    <=  16'h03C0;
                char18[11]    <=  16'h03C0;
                char18[12]    <=  16'h03C0;
                char18[13]    <=  16'h03C0;
                char18[14]    <=  16'h03C0;
                char18[15]    <=  16'h03C0;
                char18[16]    <=  16'h03C0;
                char18[17]    <=  16'h03C0;
                char18[18]    <=  16'h03C0;
                char18[19]    <=  16'h03E0;
                char18[20]    <=  16'h1FFC;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end
            4'd2  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h07E0;
                char18[5]     <=  16'h1EF8;
                char18[6]     <=  16'h383C;
                char18[7]     <=  16'h781C;
                char18[8]     <=  16'h7C1C;
                char18[9]     <=  16'h381C;
                char18[10]    <=  16'h003C;
                char18[11]    <=  16'h0038;
                char18[12]    <=  16'h0070;
                char18[13]    <=  16'h01E0;
                char18[14]    <=  16'h0380;
                char18[15]    <=  16'h0700;
                char18[16]    <=  16'h0E06;
                char18[17]    <=  16'h1C0E;
                char18[18]    <=  16'h301C;
                char18[19]    <=  16'h7FFC;
                char18[20]    <=  16'h7FFC;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h07E0;
                char18[5]     <=  16'h1EF0;
                char18[6]     <=  16'h3838;
                char18[7]     <=  16'h383C;
                char18[8]     <=  16'h383C;
                char18[9]     <=  16'h003C;
                char18[10]    <=  16'h0078;
                char18[11]    <=  16'h03F0;
                char18[12]    <=  16'h03F0;
                char18[13]    <=  16'h0038;
                char18[14]    <=  16'h001C;
                char18[15]    <=  16'h001E;
                char18[16]    <=  16'h381E;
                char18[17]    <=  16'h781E;
                char18[18]    <=  16'h783C;
                char18[19]    <=  16'h3C78;
                char18[20]    <=  16'h0FE0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h0070;
                char18[5]     <=  16'h0070;
                char18[6]     <=  16'h00F0;
                char18[7]     <=  16'h01F0;
                char18[8]     <=  16'h03F0;
                char18[9]     <=  16'h0770;
                char18[10]    <=  16'h0E70;
                char18[11]    <=  16'h0C70;
                char18[12]    <=  16'h1870;
                char18[13]    <=  16'h3070;
                char18[14]    <=  16'h7070;
                char18[15]    <=  16'hFFFF;
                char18[16]    <=  16'h0070;
                char18[17]    <=  16'h0070;
                char18[18]    <=  16'h0070;
                char18[19]    <=  16'h00F8;
                char18[20]    <=  16'h07FE;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h1FFC;
                char18[5]     <=  16'h1FFC;
                char18[6]     <=  16'h3800;
                char18[7]     <=  16'h3800;
                char18[8]     <=  16'h3800;
                char18[9]     <=  16'h3800;
                char18[10]    <=  16'h3FF0;
                char18[11]    <=  16'h3FF8;
                char18[12]    <=  16'h383C;
                char18[13]    <=  16'h101C;
                char18[14]    <=  16'h001E;
                char18[15]    <=  16'h001E;
                char18[16]    <=  16'h381E;
                char18[17]    <=  16'h781C;
                char18[18]    <=  16'h783C;
                char18[19]    <=  16'h3C78;
                char18[20]    <=  16'h0FF0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h03F0;
                char18[5]     <=  16'h0F38;
                char18[6]     <=  16'h1C3C;
                char18[7]     <=  16'h383C;
                char18[8]     <=  16'h3800;
                char18[9]     <=  16'h7800;
                char18[10]    <=  16'h7BF0;
                char18[11]    <=  16'h7FF8;
                char18[12]    <=  16'h7C3C;
                char18[13]    <=  16'h781E;
                char18[14]    <=  16'h781E;
                char18[15]    <=  16'h781E;
                char18[16]    <=  16'h781E;
                char18[17]    <=  16'h381E;
                char18[18]    <=  16'h3C1C;
                char18[19]    <=  16'h1E38;
                char18[20]    <=  16'h07F0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h3FFE;
                char18[5]     <=  16'h3FFE;
                char18[6]     <=  16'h381C;
                char18[7]     <=  16'h7018;
                char18[8]     <=  16'h7030;
                char18[9]     <=  16'h0070;
                char18[10]    <=  16'h00E0;
                char18[11]    <=  16'h00E0;
                char18[12]    <=  16'h01C0;
                char18[13]    <=  16'h01C0;
                char18[14]    <=  16'h0380;
                char18[15]    <=  16'h0380;
                char18[16]    <=  16'h0780;
                char18[17]    <=  16'h0780;
                char18[18]    <=  16'h0780;
                char18[19]    <=  16'h0780;
                char18[20]    <=  16'h0780;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h07E0;
                char18[5]     <=  16'h1E78;
                char18[6]     <=  16'h381C;
                char18[7]     <=  16'h701E;
                char18[8]     <=  16'h701E;
                char18[9]     <=  16'h781C;
                char18[10]    <=  16'h3E3C;
                char18[11]    <=  16'h1FF0;
                char18[12]    <=  16'h1FF0;
                char18[13]    <=  16'h3CF8;
                char18[14]    <=  16'h783C;
                char18[15]    <=  16'h701E;
                char18[16]    <=  16'h701E;
                char18[17]    <=  16'h701E;
                char18[18]    <=  16'h701C;
                char18[19]    <=  16'h3C38;
                char18[20]    <=  16'h0FF0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h0FE0;
                char18[5]     <=  16'h1EF8;
                char18[6]     <=  16'h3838;
                char18[7]     <=  16'h781C;
                char18[8]     <=  16'h701E;
                char18[9]     <=  16'h701E;
                char18[10]    <=  16'h701E;
                char18[11]    <=  16'h781E;
                char18[12]    <=  16'h783E;
                char18[13]    <=  16'h3FFE;
                char18[14]    <=  16'h0FDE;
                char18[15]    <=  16'h001C;
                char18[16]    <=  16'h003C;
                char18[17]    <=  16'h1838;
                char18[18]    <=  16'h3C78;
                char18[19]    <=  16'h3CF0;
                char18[20]    <=  16'h1FC0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end   
            default:begin
                char18[0]     <=  16'h0000;
                char18[1]     <=  16'h0000;
                char18[2]     <=  16'h0000;
                char18[3]     <=  16'h0000;
                char18[4]     <=  16'h07E0;
                char18[5]     <=  16'h0FF0;
                char18[6]     <=  16'h1C38;
                char18[7]     <=  16'h3C3C;
                char18[8]     <=  16'h781C;
                char18[9]     <=  16'h781E;
                char18[10]    <=  16'h781E;
                char18[11]    <=  16'h781E;
                char18[12]    <=  16'h781E;
                char18[13]    <=  16'h781E;
                char18[14]    <=  16'h781E;
                char18[15]    <=  16'h781E;
                char18[16]    <=  16'h781E;
                char18[17]    <=  16'h383C;
                char18[18]    <=  16'h3C38;
                char18[19]    <=  16'h1E78;
                char18[20]    <=  16'h07E0;
                char18[21]    <=  16'h0000;
                char18[22]    <=  16'h0000;
                char18[23]    <=  16'h0000;
            end
        endcase
//------------------------------------------------------------------------------
//--------------------------------------ppm-------------------------------------
//------------------------------------------------------------------------------
always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char24[0]     <=  16'h0000;
       char24[1]     <=  16'h0000;
       char24[2]     <=  16'h0000;
       char24[3]     <=  16'h0000;
       char24[4]     <=  16'h07E0;
       char24[5]     <=  16'h0FF0;
       char24[6]     <=  16'h1C38;
       char24[7]     <=  16'h3C3C;
       char24[8]     <=  16'h781C;
       char24[9]     <=  16'h781E;
       char24[10]    <=  16'h781E;
       char24[11]    <=  16'h781E;
       char24[12]    <=  16'h781E;
       char24[13]    <=  16'h781E;
       char24[14]    <=  16'h781E;
       char24[15]    <=  16'h781E;
       char24[16]    <=  16'h781E;
       char24[17]    <=  16'h383C;
       char24[18]    <=  16'h3C38;
       char24[19]    <=  16'h1E78;
       char24[20]    <=  16'h07E0;
       char24[21]    <=  16'h0000;
       char24[22]    <=  16'h0000;
       char24[23]    <=  16'h0000;
    end
    else    
        case(hun5)
            4'd0  :  begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h07E0;
                char24[5]     <=  16'h0FF0;
                char24[6]     <=  16'h1C38;
                char24[7]     <=  16'h3C3C;
                char24[8]     <=  16'h781C;
                char24[9]     <=  16'h781E;
                char24[10]    <=  16'h781E;
                char24[11]    <=  16'h781E;
                char24[12]    <=  16'h781E;
                char24[13]    <=  16'h781E;
                char24[14]    <=  16'h781E;
                char24[15]    <=  16'h781E;
                char24[16]    <=  16'h781E;
                char24[17]    <=  16'h383C;
                char24[18]    <=  16'h3C38;
                char24[19]    <=  16'h1E78;
                char24[20]    <=  16'h07E0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h00C0;
                char24[5]     <=  16'h0FC0;
                char24[6]     <=  16'h1FC0;
                char24[7]     <=  16'h03C0;
                char24[8]     <=  16'h03C0;
                char24[9]     <=  16'h03C0;
                char24[10]    <=  16'h03C0;
                char24[11]    <=  16'h03C0;
                char24[12]    <=  16'h03C0;
                char24[13]    <=  16'h03C0;
                char24[14]    <=  16'h03C0;
                char24[15]    <=  16'h03C0;
                char24[16]    <=  16'h03C0;
                char24[17]    <=  16'h03C0;
                char24[18]    <=  16'h03C0;
                char24[19]    <=  16'h03E0;
                char24[20]    <=  16'h1FFC;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end
            4'd2  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h07E0;
                char24[5]     <=  16'h1EF8;
                char24[6]     <=  16'h383C;
                char24[7]     <=  16'h781C;
                char24[8]     <=  16'h7C1C;
                char24[9]     <=  16'h381C;
                char24[10]    <=  16'h003C;
                char24[11]    <=  16'h0038;
                char24[12]    <=  16'h0070;
                char24[13]    <=  16'h01E0;
                char24[14]    <=  16'h0380;
                char24[15]    <=  16'h0700;
                char24[16]    <=  16'h0E06;
                char24[17]    <=  16'h1C0E;
                char24[18]    <=  16'h301C;
                char24[19]    <=  16'h7FFC;
                char24[20]    <=  16'h7FFC;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h07E0;
                char24[5]     <=  16'h1EF0;
                char24[6]     <=  16'h3838;
                char24[7]     <=  16'h383C;
                char24[8]     <=  16'h383C;
                char24[9]     <=  16'h003C;
                char24[10]    <=  16'h0078;
                char24[11]    <=  16'h03F0;
                char24[12]    <=  16'h03F0;
                char24[13]    <=  16'h0038;
                char24[14]    <=  16'h001C;
                char24[15]    <=  16'h001E;
                char24[16]    <=  16'h381E;
                char24[17]    <=  16'h781E;
                char24[18]    <=  16'h783C;
                char24[19]    <=  16'h3C78;
                char24[20]    <=  16'h0FE0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h0070;
                char24[5]     <=  16'h0070;
                char24[6]     <=  16'h00F0;
                char24[7]     <=  16'h01F0;
                char24[8]     <=  16'h03F0;
                char24[9]     <=  16'h0770;
                char24[10]    <=  16'h0E70;
                char24[11]    <=  16'h0C70;
                char24[12]    <=  16'h1870;
                char24[13]    <=  16'h3070;
                char24[14]    <=  16'h7070;
                char24[15]    <=  16'hFFFF;
                char24[16]    <=  16'h0070;
                char24[17]    <=  16'h0070;
                char24[18]    <=  16'h0070;
                char24[19]    <=  16'h00F8;
                char24[20]    <=  16'h07FE;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h1FFC;
                char24[5]     <=  16'h1FFC;
                char24[6]     <=  16'h3800;
                char24[7]     <=  16'h3800;
                char24[8]     <=  16'h3800;
                char24[9]     <=  16'h3800;
                char24[10]    <=  16'h3FF0;
                char24[11]    <=  16'h3FF8;
                char24[12]    <=  16'h383C;
                char24[13]    <=  16'h101C;
                char24[14]    <=  16'h001E;
                char24[15]    <=  16'h001E;
                char24[16]    <=  16'h381E;
                char24[17]    <=  16'h781C;
                char24[18]    <=  16'h783C;
                char24[19]    <=  16'h3C78;
                char24[20]    <=  16'h0FF0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h03F0;
                char24[5]     <=  16'h0F38;
                char24[6]     <=  16'h1C3C;
                char24[7]     <=  16'h383C;
                char24[8]     <=  16'h3800;
                char24[9]     <=  16'h7800;
                char24[10]    <=  16'h7BF0;
                char24[11]    <=  16'h7FF8;
                char24[12]    <=  16'h7C3C;
                char24[13]    <=  16'h781E;
                char24[14]    <=  16'h781E;
                char24[15]    <=  16'h781E;
                char24[16]    <=  16'h781E;
                char24[17]    <=  16'h381E;
                char24[18]    <=  16'h3C1C;
                char24[19]    <=  16'h1E38;
                char24[20]    <=  16'h07F0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h3FFE;
                char24[5]     <=  16'h3FFE;
                char24[6]     <=  16'h381C;
                char24[7]     <=  16'h7018;
                char24[8]     <=  16'h7030;
                char24[9]     <=  16'h0070;
                char24[10]    <=  16'h00E0;
                char24[11]    <=  16'h00E0;
                char24[12]    <=  16'h01C0;
                char24[13]    <=  16'h01C0;
                char24[14]    <=  16'h0380;
                char24[15]    <=  16'h0380;
                char24[16]    <=  16'h0780;
                char24[17]    <=  16'h0780;
                char24[18]    <=  16'h0780;
                char24[19]    <=  16'h0780;
                char24[20]    <=  16'h0780;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h07E0;
                char24[5]     <=  16'h1E78;
                char24[6]     <=  16'h381C;
                char24[7]     <=  16'h701E;
                char24[8]     <=  16'h701E;
                char24[9]     <=  16'h781C;
                char24[10]    <=  16'h3E3C;
                char24[11]    <=  16'h1FF0;
                char24[12]    <=  16'h1FF0;
                char24[13]    <=  16'h3CF8;
                char24[14]    <=  16'h783C;
                char24[15]    <=  16'h701E;
                char24[16]    <=  16'h701E;
                char24[17]    <=  16'h701E;
                char24[18]    <=  16'h701C;
                char24[19]    <=  16'h3C38;
                char24[20]    <=  16'h0FF0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h0FE0;
                char24[5]     <=  16'h1EF8;
                char24[6]     <=  16'h3838;
                char24[7]     <=  16'h781C;
                char24[8]     <=  16'h701E;
                char24[9]     <=  16'h701E;
                char24[10]    <=  16'h701E;
                char24[11]    <=  16'h781E;
                char24[12]    <=  16'h783E;
                char24[13]    <=  16'h3FFE;
                char24[14]    <=  16'h0FDE;
                char24[15]    <=  16'h001C;
                char24[16]    <=  16'h003C;
                char24[17]    <=  16'h1838;
                char24[18]    <=  16'h3C78;
                char24[19]    <=  16'h3CF0;
                char24[20]    <=  16'h1FC0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end   
            default:begin
                char24[0]     <=  16'h0000;
                char24[1]     <=  16'h0000;
                char24[2]     <=  16'h0000;
                char24[3]     <=  16'h0000;
                char24[4]     <=  16'h07E0;
                char24[5]     <=  16'h0FF0;
                char24[6]     <=  16'h1C38;
                char24[7]     <=  16'h3C3C;
                char24[8]     <=  16'h781C;
                char24[9]     <=  16'h781E;
                char24[10]    <=  16'h781E;
                char24[11]    <=  16'h781E;
                char24[12]    <=  16'h781E;
                char24[13]    <=  16'h781E;
                char24[14]    <=  16'h781E;
                char24[15]    <=  16'h781E;
                char24[16]    <=  16'h781E;
                char24[17]    <=  16'h383C;
                char24[18]    <=  16'h3C38;
                char24[19]    <=  16'h1E78;
                char24[20]    <=  16'h07E0;
                char24[21]    <=  16'h0000;
                char24[22]    <=  16'h0000;
                char24[23]    <=  16'h0000;
            end
        endcase
always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char25[0]     <=  16'h0000;
       char25[1]     <=  16'h0000;
       char25[2]     <=  16'h0000;
       char25[3]     <=  16'h0000;
       char25[4]     <=  16'h07E0;
       char25[5]     <=  16'h0FF0;
       char25[6]     <=  16'h1C38;
       char25[7]     <=  16'h3C3C;
       char25[8]     <=  16'h781C;
       char25[9]     <=  16'h781E;
       char25[10]    <=  16'h781E;
       char25[11]    <=  16'h781E;
       char25[12]    <=  16'h781E;
       char25[13]    <=  16'h781E;
       char25[14]    <=  16'h781E;
       char25[15]    <=  16'h781E;
       char25[16]    <=  16'h781E;
       char25[17]    <=  16'h383C;
       char25[18]    <=  16'h3C38;
       char25[19]    <=  16'h1E78;
       char25[20]    <=  16'h07E0;
       char25[21]    <=  16'h0000;
       char25[22]    <=  16'h0000;
       char25[23]    <=  16'h0000;
    end
    else    
        case(ten5)
            4'd0  :  begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h07E0;
                char25[5]     <=  16'h0FF0;
                char25[6]     <=  16'h1C38;
                char25[7]     <=  16'h3C3C;
                char25[8]     <=  16'h781C;
                char25[9]     <=  16'h781E;
                char25[10]    <=  16'h781E;
                char25[11]    <=  16'h781E;
                char25[12]    <=  16'h781E;
                char25[13]    <=  16'h781E;
                char25[14]    <=  16'h781E;
                char25[15]    <=  16'h781E;
                char25[16]    <=  16'h781E;
                char25[17]    <=  16'h383C;
                char25[18]    <=  16'h3C38;
                char25[19]    <=  16'h1E78;
                char25[20]    <=  16'h07E0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h00C0;
                char25[5]     <=  16'h0FC0;
                char25[6]     <=  16'h1FC0;
                char25[7]     <=  16'h03C0;
                char25[8]     <=  16'h03C0;
                char25[9]     <=  16'h03C0;
                char25[10]    <=  16'h03C0;
                char25[11]    <=  16'h03C0;
                char25[12]    <=  16'h03C0;
                char25[13]    <=  16'h03C0;
                char25[14]    <=  16'h03C0;
                char25[15]    <=  16'h03C0;
                char25[16]    <=  16'h03C0;
                char25[17]    <=  16'h03C0;
                char25[18]    <=  16'h03C0;
                char25[19]    <=  16'h03E0;
                char25[20]    <=  16'h1FFC;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end
            4'd2  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h07E0;
                char25[5]     <=  16'h1EF8;
                char25[6]     <=  16'h383C;
                char25[7]     <=  16'h781C;
                char25[8]     <=  16'h7C1C;
                char25[9]     <=  16'h381C;
                char25[10]    <=  16'h003C;
                char25[11]    <=  16'h0038;
                char25[12]    <=  16'h0070;
                char25[13]    <=  16'h01E0;
                char25[14]    <=  16'h0380;
                char25[15]    <=  16'h0700;
                char25[16]    <=  16'h0E06;
                char25[17]    <=  16'h1C0E;
                char25[18]    <=  16'h301C;
                char25[19]    <=  16'h7FFC;
                char25[20]    <=  16'h7FFC;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h07E0;
                char25[5]     <=  16'h1EF0;
                char25[6]     <=  16'h3838;
                char25[7]     <=  16'h383C;
                char25[8]     <=  16'h383C;
                char25[9]     <=  16'h003C;
                char25[10]    <=  16'h0078;
                char25[11]    <=  16'h03F0;
                char25[12]    <=  16'h03F0;
                char25[13]    <=  16'h0038;
                char25[14]    <=  16'h001C;
                char25[15]    <=  16'h001E;
                char25[16]    <=  16'h381E;
                char25[17]    <=  16'h781E;
                char25[18]    <=  16'h783C;
                char25[19]    <=  16'h3C78;
                char25[20]    <=  16'h0FE0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h0070;
                char25[5]     <=  16'h0070;
                char25[6]     <=  16'h00F0;
                char25[7]     <=  16'h01F0;
                char25[8]     <=  16'h03F0;
                char25[9]     <=  16'h0770;
                char25[10]    <=  16'h0E70;
                char25[11]    <=  16'h0C70;
                char25[12]    <=  16'h1870;
                char25[13]    <=  16'h3070;
                char25[14]    <=  16'h7070;
                char25[15]    <=  16'hFFFF;
                char25[16]    <=  16'h0070;
                char25[17]    <=  16'h0070;
                char25[18]    <=  16'h0070;
                char25[19]    <=  16'h00F8;
                char25[20]    <=  16'h07FE;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h1FFC;
                char25[5]     <=  16'h1FFC;
                char25[6]     <=  16'h3800;
                char25[7]     <=  16'h3800;
                char25[8]     <=  16'h3800;
                char25[9]     <=  16'h3800;
                char25[10]    <=  16'h3FF0;
                char25[11]    <=  16'h3FF8;
                char25[12]    <=  16'h383C;
                char25[13]    <=  16'h101C;
                char25[14]    <=  16'h001E;
                char25[15]    <=  16'h001E;
                char25[16]    <=  16'h381E;
                char25[17]    <=  16'h781C;
                char25[18]    <=  16'h783C;
                char25[19]    <=  16'h3C78;
                char25[20]    <=  16'h0FF0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h03F0;
                char25[5]     <=  16'h0F38;
                char25[6]     <=  16'h1C3C;
                char25[7]     <=  16'h383C;
                char25[8]     <=  16'h3800;
                char25[9]     <=  16'h7800;
                char25[10]    <=  16'h7BF0;
                char25[11]    <=  16'h7FF8;
                char25[12]    <=  16'h7C3C;
                char25[13]    <=  16'h781E;
                char25[14]    <=  16'h781E;
                char25[15]    <=  16'h781E;
                char25[16]    <=  16'h781E;
                char25[17]    <=  16'h381E;
                char25[18]    <=  16'h3C1C;
                char25[19]    <=  16'h1E38;
                char25[20]    <=  16'h07F0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h3FFE;
                char25[5]     <=  16'h3FFE;
                char25[6]     <=  16'h381C;
                char25[7]     <=  16'h7018;
                char25[8]     <=  16'h7030;
                char25[9]     <=  16'h0070;
                char25[10]    <=  16'h00E0;
                char25[11]    <=  16'h00E0;
                char25[12]    <=  16'h01C0;
                char25[13]    <=  16'h01C0;
                char25[14]    <=  16'h0380;
                char25[15]    <=  16'h0380;
                char25[16]    <=  16'h0780;
                char25[17]    <=  16'h0780;
                char25[18]    <=  16'h0780;
                char25[19]    <=  16'h0780;
                char25[20]    <=  16'h0780;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h07E0;
                char25[5]     <=  16'h1E78;
                char25[6]     <=  16'h381C;
                char25[7]     <=  16'h701E;
                char25[8]     <=  16'h701E;
                char25[9]     <=  16'h781C;
                char25[10]    <=  16'h3E3C;
                char25[11]    <=  16'h1FF0;
                char25[12]    <=  16'h1FF0;
                char25[13]    <=  16'h3CF8;
                char25[14]    <=  16'h783C;
                char25[15]    <=  16'h701E;
                char25[16]    <=  16'h701E;
                char25[17]    <=  16'h701E;
                char25[18]    <=  16'h701C;
                char25[19]    <=  16'h3C38;
                char25[20]    <=  16'h0FF0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h0FE0;
                char25[5]     <=  16'h1EF8;
                char25[6]     <=  16'h3838;
                char25[7]     <=  16'h781C;
                char25[8]     <=  16'h701E;
                char25[9]     <=  16'h701E;
                char25[10]    <=  16'h701E;
                char25[11]    <=  16'h781E;
                char25[12]    <=  16'h783E;
                char25[13]    <=  16'h3FFE;
                char25[14]    <=  16'h0FDE;
                char25[15]    <=  16'h001C;
                char25[16]    <=  16'h003C;
                char25[17]    <=  16'h1838;
                char25[18]    <=  16'h3C78;
                char25[19]    <=  16'h3CF0;
                char25[20]    <=  16'h1FC0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end   
            default:begin
                char25[0]     <=  16'h0000;
                char25[1]     <=  16'h0000;
                char25[2]     <=  16'h0000;
                char25[3]     <=  16'h0000;
                char25[4]     <=  16'h07E0;
                char25[5]     <=  16'h0FF0;
                char25[6]     <=  16'h1C38;
                char25[7]     <=  16'h3C3C;
                char25[8]     <=  16'h781C;
                char25[9]     <=  16'h781E;
                char25[10]    <=  16'h781E;
                char25[11]    <=  16'h781E;
                char25[12]    <=  16'h781E;
                char25[13]    <=  16'h781E;
                char25[14]    <=  16'h781E;
                char25[15]    <=  16'h781E;
                char25[16]    <=  16'h781E;
                char25[17]    <=  16'h383C;
                char25[18]    <=  16'h3C38;
                char25[19]    <=  16'h1E78;
                char25[20]    <=  16'h07E0;
                char25[21]    <=  16'h0000;
                char25[22]    <=  16'h0000;
                char25[23]    <=  16'h0000;
            end
        endcase

always@(posedge tft_clk_33m or  negedge sys_rst_n)
    if(!sys_rst_n)begin
       char26[0]     <=  16'h0000;
       char26[1]     <=  16'h0000;
       char26[2]     <=  16'h0000;
       char26[3]     <=  16'h0000;
       char26[4]     <=  16'h07E0;
       char26[5]     <=  16'h0FF0;
       char26[6]     <=  16'h1C38;
       char26[7]     <=  16'h3C3C;
       char26[8]     <=  16'h781C;
       char26[9]     <=  16'h781E;
       char26[10]    <=  16'h781E;
       char26[11]    <=  16'h781E;
       char26[12]    <=  16'h781E;
       char26[13]    <=  16'h781E;
       char26[14]    <=  16'h781E;
       char26[15]    <=  16'h781E;
       char26[16]    <=  16'h781E;
       char26[17]    <=  16'h383C;
       char26[18]    <=  16'h3C38;
       char26[19]    <=  16'h1E78;
       char26[20]    <=  16'h07E0;
       char26[21]    <=  16'h0000;
       char26[22]    <=  16'h0000;
       char26[23]    <=  16'h0000;
    end
    else    
        case(unit5)
            4'd0  :  begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h07E0;
                char26[5]     <=  16'h0FF0;
                char26[6]     <=  16'h1C38;
                char26[7]     <=  16'h3C3C;
                char26[8]     <=  16'h781C;
                char26[9]     <=  16'h781E;
                char26[10]    <=  16'h781E;
                char26[11]    <=  16'h781E;
                char26[12]    <=  16'h781E;
                char26[13]    <=  16'h781E;
                char26[14]    <=  16'h781E;
                char26[15]    <=  16'h781E;
                char26[16]    <=  16'h781E;
                char26[17]    <=  16'h383C;
                char26[18]    <=  16'h3C38;
                char26[19]    <=  16'h1E78;
                char26[20]    <=  16'h07E0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
                end
            4'd1  :  begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h00C0;
                char26[5]     <=  16'h0FC0;
                char26[6]     <=  16'h1FC0;
                char26[7]     <=  16'h03C0;
                char26[8]     <=  16'h03C0;
                char26[9]     <=  16'h03C0;
                char26[10]    <=  16'h03C0;
                char26[11]    <=  16'h03C0;
                char26[12]    <=  16'h03C0;
                char26[13]    <=  16'h03C0;
                char26[14]    <=  16'h03C0;
                char26[15]    <=  16'h03C0;
                char26[16]    <=  16'h03C0;
                char26[17]    <=  16'h03C0;
                char26[18]    <=  16'h03C0;
                char26[19]    <=  16'h03E0;
                char26[20]    <=  16'h1FFC;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end
            4'd2  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h07E0;
                char26[5]     <=  16'h1EF8;
                char26[6]     <=  16'h383C;
                char26[7]     <=  16'h781C;
                char26[8]     <=  16'h7C1C;
                char26[9]     <=  16'h381C;
                char26[10]    <=  16'h003C;
                char26[11]    <=  16'h0038;
                char26[12]    <=  16'h0070;
                char26[13]    <=  16'h01E0;
                char26[14]    <=  16'h0380;
                char26[15]    <=  16'h0700;
                char26[16]    <=  16'h0E06;
                char26[17]    <=  16'h1C0E;
                char26[18]    <=  16'h301C;
                char26[19]    <=  16'h7FFC;
                char26[20]    <=  16'h7FFC;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end 
            4'd3  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h07E0;
                char26[5]     <=  16'h1EF0;
                char26[6]     <=  16'h3838;
                char26[7]     <=  16'h383C;
                char26[8]     <=  16'h383C;
                char26[9]     <=  16'h003C;
                char26[10]    <=  16'h0078;
                char26[11]    <=  16'h03F0;
                char26[12]    <=  16'h03F0;
                char26[13]    <=  16'h0038;
                char26[14]    <=  16'h001C;
                char26[15]    <=  16'h001E;
                char26[16]    <=  16'h381E;
                char26[17]    <=  16'h781E;
                char26[18]    <=  16'h783C;
                char26[19]    <=  16'h3C78;
                char26[20]    <=  16'h0FE0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end   
            4'd4  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h0070;
                char26[5]     <=  16'h0070;
                char26[6]     <=  16'h00F0;
                char26[7]     <=  16'h01F0;
                char26[8]     <=  16'h03F0;
                char26[9]     <=  16'h0770;
                char26[10]    <=  16'h0E70;
                char26[11]    <=  16'h0C70;
                char26[12]    <=  16'h1870;
                char26[13]    <=  16'h3070;
                char26[14]    <=  16'h7070;
                char26[15]    <=  16'hFFFF;
                char26[16]    <=  16'h0070;
                char26[17]    <=  16'h0070;
                char26[18]    <=  16'h0070;
                char26[19]    <=  16'h00F8;
                char26[20]    <=  16'h07FE;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end   
            4'd5  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h1FFC;
                char26[5]     <=  16'h1FFC;
                char26[6]     <=  16'h3800;
                char26[7]     <=  16'h3800;
                char26[8]     <=  16'h3800;
                char26[9]     <=  16'h3800;
                char26[10]    <=  16'h3FF0;
                char26[11]    <=  16'h3FF8;
                char26[12]    <=  16'h383C;
                char26[13]    <=  16'h101C;
                char26[14]    <=  16'h001E;
                char26[15]    <=  16'h001E;
                char26[16]    <=  16'h381E;
                char26[17]    <=  16'h781C;
                char26[18]    <=  16'h783C;
                char26[19]    <=  16'h3C78;
                char26[20]    <=  16'h0FF0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end   
            4'd6  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h03F0;
                char26[5]     <=  16'h0F38;
                char26[6]     <=  16'h1C3C;
                char26[7]     <=  16'h383C;
                char26[8]     <=  16'h3800;
                char26[9]     <=  16'h7800;
                char26[10]    <=  16'h7BF0;
                char26[11]    <=  16'h7FF8;
                char26[12]    <=  16'h7C3C;
                char26[13]    <=  16'h781E;
                char26[14]    <=  16'h781E;
                char26[15]    <=  16'h781E;
                char26[16]    <=  16'h781E;
                char26[17]    <=  16'h381E;
                char26[18]    <=  16'h3C1C;
                char26[19]    <=  16'h1E38;
                char26[20]    <=  16'h07F0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;               
            end   
            4'd7  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h3FFE;
                char26[5]     <=  16'h3FFE;
                char26[6]     <=  16'h381C;
                char26[7]     <=  16'h7018;
                char26[8]     <=  16'h7030;
                char26[9]     <=  16'h0070;
                char26[10]    <=  16'h00E0;
                char26[11]    <=  16'h00E0;
                char26[12]    <=  16'h01C0;
                char26[13]    <=  16'h01C0;
                char26[14]    <=  16'h0380;
                char26[15]    <=  16'h0380;
                char26[16]    <=  16'h0780;
                char26[17]    <=  16'h0780;
                char26[18]    <=  16'h0780;
                char26[19]    <=  16'h0780;
                char26[20]    <=  16'h0780;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end   
            4'd8  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h07E0;
                char26[5]     <=  16'h1E78;
                char26[6]     <=  16'h381C;
                char26[7]     <=  16'h701E;
                char26[8]     <=  16'h701E;
                char26[9]     <=  16'h781C;
                char26[10]    <=  16'h3E3C;
                char26[11]    <=  16'h1FF0;
                char26[12]    <=  16'h1FF0;
                char26[13]    <=  16'h3CF8;
                char26[14]    <=  16'h783C;
                char26[15]    <=  16'h701E;
                char26[16]    <=  16'h701E;
                char26[17]    <=  16'h701E;
                char26[18]    <=  16'h701C;
                char26[19]    <=  16'h3C38;
                char26[20]    <=  16'h0FF0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end   
            4'd9  : begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h0FE0;
                char26[5]     <=  16'h1EF8;
                char26[6]     <=  16'h3838;
                char26[7]     <=  16'h781C;
                char26[8]     <=  16'h701E;
                char26[9]     <=  16'h701E;
                char26[10]    <=  16'h701E;
                char26[11]    <=  16'h781E;
                char26[12]    <=  16'h783E;
                char26[13]    <=  16'h3FFE;
                char26[14]    <=  16'h0FDE;
                char26[15]    <=  16'h001C;
                char26[16]    <=  16'h003C;
                char26[17]    <=  16'h1838;
                char26[18]    <=  16'h3C78;
                char26[19]    <=  16'h3CF0;
                char26[20]    <=  16'h1FC0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end   
            default:begin
                char26[0]     <=  16'h0000;
                char26[1]     <=  16'h0000;
                char26[2]     <=  16'h0000;
                char26[3]     <=  16'h0000;
                char26[4]     <=  16'h07E0;
                char26[5]     <=  16'h0FF0;
                char26[6]     <=  16'h1C38;
                char26[7]     <=  16'h3C3C;
                char26[8]     <=  16'h781C;
                char26[9]     <=  16'h781E;
                char26[10]    <=  16'h781E;
                char26[11]    <=  16'h781E;
                char26[12]    <=  16'h781E;
                char26[13]    <=  16'h781E;
                char26[14]    <=  16'h781E;
                char26[15]    <=  16'h781E;
                char26[16]    <=  16'h781E;
                char26[17]    <=  16'h383C;
                char26[18]    <=  16'h3C38;
                char26[19]    <=  16'h1E78;
                char26[20]    <=  16'h07E0;
                char26[21]    <=  16'h0000;
                char26[22]    <=  16'h0000;
                char26[23]    <=  16'h0000;
            end
        endcase
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
//-----------------------------------AD图像显示----------------------------------
//------------------------------------------------------------------------------
parameter CNT_MAX = 26'd66_666_664;

reg [25:0] cnt ;
reg cnt_flag ;
reg [9:0] charx ;

always@(posedge tft_clk_33m or negedge sys_rst_n)begin
    if(!sys_rst_n)
        cnt   <= 25'd0;
    else if(cnt == CNT_MAX)
        cnt <= 25'b0;
    else
        cnt <= cnt + 1'b1;
end

 always@(posedge tft_clk_33m or negedge sys_rst_n)begin
    if(!sys_rst_n)
        cnt_flag <= 1'b0;
    else if(cnt == CNT_MAX - 3)
        cnt_flag <= 1'b1;
    else
        cnt_flag <= 1'b0;
 end


 always@(posedge tft_clk_33m or negedge sys_rst_n)begin
    if(!sys_rst_n)
        charx <= 10'd0;
    else if(charx == 10'd720 && cnt_flag == 1'b1)
        charx <= 10'd0;
    else if(cnt_flag == 1'b1)
        charx <= charx +10'd1;
    else
        charx <= charx;
 end

// assign rdaddress =pix_x+(pix_y-10'd32)*800;
// assign wraddress =charx+(10'd384-ch1)*800;
reg [18:0]rdaddress;
reg [18:0]wraddress;
always@(posedge tft_clk_33m or negedge sys_rst_n)begin
   if(!sys_rst_n) begin
       rdaddress <=0;
       wraddress <=0;
   end
   else begin
       rdaddress <=pix_x-10'd50+(pix_y-10'd30)*720;
       wraddress <=charx+(10'd340-data_out)*720;
   end
   end


ram9	ram9_inst (
	.clock ( tft_clk_33m ),
	.data ( 1'b1 ),
	.rdaddress ( rdaddress ),
	.rden ( 1 ),
	.wraddress ( wraddress ),
	.wren ( 1 ),
	.q ( q )
	);

parameter CNT_MAX1 = 27'd133_333_332;

reg [26:0] cnt1 ;
reg cnt_flag1 ;
reg [8:0] charx1 ;

always@(posedge tft_clk_33m or negedge sys_rst_n)begin
    if(!sys_rst_n)
        cnt1   <= 25'd0;
    else if(cnt == CNT_MAX1)
        cnt1 <= 25'b0;
    else
        cnt1 <= cnt1 + 1'b1;
end

 always@(posedge tft_clk_33m or negedge sys_rst_n)begin
    if(!sys_rst_n)
        cnt_flag1 <= 1'b0;
    else if(cnt1 == CNT_MAX1 - 3)
        cnt_flag1 <= 1'b1;
    else
        cnt_flag1 <= 1'b0;
 end


 always@(posedge tft_clk_33m or negedge sys_rst_n)begin
    if(!sys_rst_n)
        charx1 <= 10'd0;
    else if(charx1 == 10'd300 && cnt_flag1 == 1'b1)
        charx1 <= 10'd0;
    else if(cnt_flag1 == 1'b1)
        charx1 <= charx1 +10'd1;
    else
        charx1 <= charx1;
 end



//ch1
reg [15:0]rdaddress1;
reg [15:0]wraddress1;
always@(posedge tft_clk_33m or negedge sys_rst_n)begin
   if(!sys_rst_n) begin
       rdaddress1 <=0;
       wraddress1 <=0;
   end
   else begin
       rdaddress1 <=pix_x-10'd50+(pix_y-10'd50)*280;
       wraddress1 <=charx1+(10'd114-(ch1>>1))*280;
   end
   end

ram1	ram1_inst (
	.clock ( tft_clk_33m ),
	.data ( 1'b1 ),
	.rdaddress ( rdaddress1 ),
	.rden ( 1 ),
	.wraddress ( wraddress1 ),
	.wren ( 1 ),
	.q ( q1 )
	);

//ch2
reg [15:0]rdaddress2;
reg [15:0]wraddress2;
always@(posedge tft_clk_33m or negedge sys_rst_n)begin
   if(!sys_rst_n) begin
       rdaddress2 <=0;
       wraddress2 <=0;
   end
   else begin
       rdaddress2 <=pix_x-10'd450+(pix_y-10'd50)*280;
       wraddress2 <=charx1+(10'd114-(ch2>>1))*280;
   end
   end

ram2	ram2_inst (
	.clock ( tft_clk_33m ),
	.data ( 1'b1 ),
	.rdaddress ( rdaddress2 ),
	.rden ( 1 ),
	.wraddress ( wraddress2 ),
	.wren ( 1 ),
	.q ( q2 )
	);

//ch3
reg [15:0]rdaddress3;
reg [15:0]wraddress3;
always@(posedge tft_clk_33m or negedge sys_rst_n)begin
   if(!sys_rst_n) begin
       rdaddress3 <=0;
       wraddress3 <=0;
   end
   else begin
       rdaddress3 <=pix_x-10'd50+(pix_y-10'd230)*280;
       wraddress3 <=charx1+(10'd114-(ch3>>1))*280;
   end
   end

ram3	ram3_inst (
	.clock ( tft_clk_33m ),
	.data ( 1'b1 ),
	.rdaddress ( rdaddress3 ),
	.rden ( 1 ),
	.wraddress ( wraddress3 ),
	.wren ( 1 ),
	.q ( q3 )
	);

//ch4
reg [15:0]rdaddress4;
reg [15:0]wraddress4;
always@(posedge tft_clk_33m or negedge sys_rst_n)begin
   if(!sys_rst_n) begin
       rdaddress4 <=0;
       wraddress4 <=0;
   end
   else begin
       rdaddress4 <=pix_x-10'd450+(pix_y-10'd230)*280;
       wraddress4 <=charx1+(10'd114-(ch4>>1))*280;
   end
   end

ram4	ram4_inst (
	.clock ( tft_clk_33m ),
	.data ( 1'b1 ),
	.rdaddress ( rdaddress4 ),
	.rden ( 1 ),
	.wraddress ( wraddress4 ),
	.wren ( 1 ),
	.q ( q4 )
	);















//--------------------------------------------------------------------------------
//-----------------------------------界面边框显示----------------------------------
//--------------------------------------------------------------------------------
// rom_font rf(
// 		.address(address),
// 		.clock(VGA_CLK/*clk_vga*/),
// 		.q(font)
// );
// wire [8:0]font;

// always @(VGA_CLK)begin
// 	 block_addr <= (v_addr >> 4) * 70 + ((h_addr) / 9);
// 	 address <= (ram_vga_ret << 4) + (v_addr % 16);

// 	 if(font[(h_addr) % 9] == 1'b1)
// 		data <= 24'hffffff;
// 	 else
// 		data <= 24'h000000;
// end	
//----------------------------------------------------------------------------------------------
//-----------------------------------pix_data:输出像素点色彩信息----------------------------------
//----------------------------------------------------------------------------------------------

always@(posedge tft_clk_33m or negedge sys_rst_n)
    if(!sys_rst_n)
        pix_data    <= BLACK;
// //JLU Gas SENSOR        
//     else    if(((pix_x >= CHAR_x1) && (pix_x < (CHAR_x1 + 10'd224)))
//                             && ((pix_y >= CHAR_y1) && (pix_y < (CHAR_y1 + 10'd24))))
//                 begin
//                     if(char1[char1_y][10'd224 - char1_x] == 1'b1)
//                         pix_data    <=  GOLDEN;
//                     else
//                         pix_data    <=  BLACK;
//                 end

//CH1
    else    if(((pix_x >= 10) && (pix_x < 10'd74))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char3[char3_y][10'd64 - char3_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH2
    else    if(((pix_x >= 10'd200) && (pix_x < (10'd264)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char19[char19_y][10'd64 - char19_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//CH3
    else    if(((pix_x >= 10'd400) && (pix_x < (10'd464)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char20[char20_y][10'd64 - char20_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end


//CH4
    else    if(((pix_x >= 10'd600) && (pix_x < (10'd664)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char21[char21_y][10'd64 - char21_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//CH1百位
    else    if(((pix_x >= 10'd74) && (pix_x < (10'd90)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char5[char5_y][10'd80 - char5_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH1十位
    else    if(((pix_x >= 10'd90) && (pix_x < (10'd106)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char6[char6_y][10'd16 - char6_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH1个位
    else    if(((pix_x >= 10'd106) && (pix_x < (10'd122)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char7[char7_y][10'd16 - char7_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//CH2百位
    else    if(((pix_x >= 10'd264) && (pix_x < (10'd280)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char10[char10_y][10'd16 - char10_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH2十位
    else    if(((pix_x >= 10'd280) && (pix_x < (10'd296)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char11[char11_y][10'd16 - char11_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH2个位
    else    if(((pix_x >= 10'd296) && (pix_x < (10'd312)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char12[char12_y][10'd16 - char12_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//CH3百位
    else    if(((pix_x >= 10'd464) && (pix_x < (10'd480)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char13[char13_y][10'd16 - char13_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH3十位
    else    if(((pix_x >= 10'd480) && (pix_x < (10'd496)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char14[char14_y][10'd16 - char14_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//CH3个位
    else    if(((pix_x >= 10'd496) && (pix_x < (10'd512)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char15[char15_y][10'd16 - char15_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//CH4百位
    else    if(((pix_x >= 10'd664) && (pix_x < (10'd680)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char16[char16_y][10'd16 - char16_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH4十位
    else    if(((pix_x >= 10'd680) && (pix_x < (10'd696)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char17[char17_y][10'd16 - char17_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//CH4个位
    else    if(((pix_x >= 10'd696) && (pix_x < (10'd712)))
                    && ((pix_y >= CHAR_y3) && (pix_y < 10'd440)))
        begin
            if(char18[char18_y][10'd16 - char18_x] == 1'b1)
                pix_data    <= WHITE;
            else
                pix_data    <=  BLACK;
        end

//ppm百位
    else    if(((pix_x >= 10'd74) && (pix_x < (10'd90)))
                    && ((pix_y >= 10'd448) && (pix_y < 10'd472)))
        begin
            if(char24[char24_y][10'd16 - char24_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//ppm十位
    else    if(((pix_x >= 10'd90) && (pix_x < (10'd106)))
                    && ((pix_y >= 10'd448) && (pix_y < 10'd472)))
        begin
            if(char25[char25_y][10'd16 - char25_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//pp,个位
    else    if(((pix_x >= 10'd106) && (pix_x < (10'd122)))
                    && ((pix_y >= 10'd448) && (pix_y < 10'd472)))
        begin
            if(char26[char26_y][10'd16 - char26_x] == 1'b1)
                pix_data    <= WHITE;
            else
                pix_data    <=  BLACK;
        end

//NH3
    else    if(((pix_x >= 10'd10) && (pix_x < ( 10'd74)))
                    && ((pix_y >= CHAR_y4) && (pix_y < 10'd472)))
        begin
            if(char4[char4_y][10'd64 - char4_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
//氨气单位
    else    if(((pix_x >= 10'd122) && (pix_x < (10'd170)))
                    && ((pix_y >= 10'd448) && (pix_y < 10'd472)))
        begin
            if(char23[char23_y][10'd48 - char23_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end


//刻度字       
    else    if (((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd71) && (pix_y < 10'd95))&& data_flag != 3'd4)
        begin
            if(char27[char27_y][10'd48 - char27_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
    else    if(((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd171) && (pix_y < 10'd195))&& data_flag != 3'd4)
        begin
            if(char28[char28_y][10'd48 - char28_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
    else    if(((pix_x >= 10'd0) && (pix_x < (10'd48)))
                    && ((pix_y >= 10'd271) && (pix_y < 10'd295))&& data_flag != 3'd4)
        begin
            if(char29[char29_y][10'd48 - char29_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
    else    if(((pix_x >= 10'd16) && (pix_x < (10'd32)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395))&& data_flag != 3'd4)
        begin
            if(char30[char30_y][10'd16 - char30_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
    else    if(((pix_x >= 10'd352) && (pix_x < (10'd448)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395))&& data_flag != 3'd4)
        begin
            if(char31[char31_y][10'd96 - char31_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end
    else    if(((pix_x >= 10'd652) && (pix_x < (10'd748)))
                    && ((pix_y >= 10'd371) && (pix_y < 10'd395))&& data_flag != 3'd4)
        begin
            if(char32[char32_y][10'd96 - char32_x] == 1'b1)
                pix_data    <=  WHITE;
            else
                pix_data    <=  BLACK;
        end

//AD图像        
    else    if(((pix_x >= 10'd50) && (pix_x < ( 10'd770)))
                && ((pix_y >= 10'd30) && (pix_y < (10'd370)))&& data_flag != 3'd4)
    begin   if (data_flag==2'd0)
	            if(q)
	    	        pix_data <= BLACK;
	            else
	    	        pix_data <= WHITE;
            else if (data_flag==2'd1)
	            if(q)
	    	        pix_data <= RED;
	            else
	    	        pix_data <= WHITE;
            else if (data_flag==2'd2)
	            if(q)
	    	        pix_data <= BLUE;
	            else
	    	        pix_data <= WHITE;
            else if (data_flag==2'd3)
	            if(q)
	    	        pix_data <= GOLDEN;
	            else
	    	        pix_data <= WHITE; 
                else
                    pix_data    <=  WHITE;       
    end
//分割线        
    else    if(pix_y==11'd400 && pix_x >= 10'd5 && pix_x < 10'd795||pix_y==11'd479 && pix_x >= 10'd5 && pix_x < 10'd795
        || pix_x==11'd5 && pix_y >= 10'd400 && pix_y < 10'd479||pix_x==11'd795 && pix_y >= 10'd400 && pix_y < 10'd479
        )
                pix_data    <=  WHITE;   

    else    if((pix_y==11'd29 && pix_x >= 10'd50 && pix_x < 10'd770||pix_y==11'd370 && pix_x >= 10'd50 && pix_x < 10'd770
        || pix_x==11'd49 && pix_y >= 10'd30 && pix_y < 10'd370||pix_x==11'd770 && pix_y >= 10'd30 && pix_y < 10'd370
        ||pix_x==11'd350 && pix_y >= 10'd371 && pix_y < 10'd380||pix_x==11'd650 && pix_y >= 10'd371 && pix_y < 10'd380
        ||pix_y==11'd70 && pix_x >= 10'd40 && pix_x < 10'd50
        ||pix_y==11'd170 && pix_x >= 10'd40 && pix_x < 10'd50
        ||pix_y==11'd270 && pix_x >= 10'd40 && pix_x < 10'd50)&& data_flag != 3'd4
        )
                pix_data    <=  WHITE;  

        


    else    if( (pix_x>=11'd5 &&pix_x<=11'd795&& pix_y >= 10'd5 && pix_y < 10'd399)&& data_flag == 3'd4) begin
            if(((pix_x >= 10'd50) && (pix_x < ( 10'd330)))
                && ((pix_y >= 10'd50) && (pix_y < (10'd164))))
	            if(q1)
	    	        pix_data <= BLACK;
	            else
	    	        pix_data <= WHITE; 

            else if(((pix_x >= 10'd450) && (pix_x < ( 10'd730)))
                && ((pix_y >= 10'd50) && (pix_y < (10'd164))))
	            if(q2)
	    	        pix_data <= RED;
	            else
	    	        pix_data <= WHITE; 

            else if(((pix_x >= 10'd50) && (pix_x < ( 10'd330)))
                && ((pix_y >= 10'd230) && (pix_y < (10'd344))))
	            if(q3)
	    	        pix_data <= BLUE;
	            else
	    	        pix_data <= WHITE; 

            else if(((pix_x >= 10'd450) && (pix_x < ( 10'd730)))
                && ((pix_y >= 10'd230) && (pix_y < (10'd344))))
	            if(q4)
	    	        pix_data <= GOLDEN;
	            else
	    	        pix_data <= WHITE;   


            else if (((pix_x >= 10'd201) && (pix_x < (10'd249)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))

                    if(char33[char33_y][10'd48 - char33_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if (((pix_x >= 10'd601) && (pix_x < (10'd649)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))

                    if(char33[char34_y][10'd48 - char34_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if (((pix_x >= 10'd201) && (pix_x < (10'd249)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))

                    if(char33[char35_y][10'd48 - char35_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if  (((pix_x >= 10'd601) && (pix_x < (10'd649)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))

                    if(char33[char36_y][10'd48 - char36_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;

            else if  (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))

                    if(char34[char37_y][10'd24 - char37_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if  (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd165) && (pix_y < 10'd181)))

                    if(char34[char38_y][10'd24 - char38_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if   (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))

                    if(char34[char39_y][10'd24 - char39_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if  (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd345) && (pix_y < 10'd361)))

                    if(char34[char40_y][10'd24 - char40_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;

            else if  (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd115) && (pix_y < 10'd131)))

                    if(char35[char41_y][10'd24 - char41_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd115) && (pix_y < 10'd131)))

                    if(char35[char42_y][10'd24 - char42_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if (((pix_x >= 10'd21) && (pix_x < (10'd45)))
                    && ((pix_y >= 10'd295) && (pix_y < 10'd311)))

                    if(char35[char43_y][10'd24 - char43_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;
            else if  (((pix_x >= 10'd421) && (pix_x < (10'd445)))
                    && ((pix_y >= 10'd295) && (pix_y < 10'd311)))

                    if(char35[char44_y][10'd24 - char44_x] == 1'b1)
                        pix_data    <=  WHITE;
                    else
                        pix_data    <=  BLACK;

            else    if(pix_x==11'd200 && pix_y >= 10'd165 && pix_y < 10'd170
                    ||pix_x==11'd200 && pix_y >= 10'd345 && pix_y < 10'd350
                    ||pix_x==11'd600 && pix_y >= 10'd165 && pix_y < 10'd170
                    ||pix_x==11'd600 && pix_y >= 10'd345 && pix_y < 10'd350

                    || pix_y==11'd114 && pix_x >= 10'd45 && pix_x < 10'd50
                    || pix_y==11'd114 && pix_x >= 10'd445 && pix_x < 10'd450
                    || pix_y==11'd294 && pix_x >= 10'd45 && pix_x < 10'd50
                    || pix_y==11'd294 && pix_x >= 10'd445 && pix_x < 10'd450
                    )
                    pix_data    <=  WHITE; 
            else
                    pix_data <= BLACK;        
    end


    else
        pix_data    <=  BLACK;

endmodule
